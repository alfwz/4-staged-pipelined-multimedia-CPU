-------------------------------------------------------------------------------
--
-- Title       : 
-- Design      : project
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- File        : F:\project345\compile\block_diagram.vhd
-- Generated   : Tue Dec  3 15:48:30 2019
-- From        : F:\project345\src\block_diagram.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_unsigned.all;

-- Included from components --
library WORK;
use work.insbuffer_type.all;

entity block_diagram is
  port(
       clk : in STD_LOGIC;
       instruction : in insBuffer(63 downto 0)
  );
end block_diagram;

architecture block_diagram of block_diagram is

---- Component declarations -----

component alu
  port (
       clk : in STD_LOGIC;
       ins : in STD_LOGIC_VECTOR(24 downto 0);
       r1 : in STD_LOGIC_VECTOR(127 downto 0);
       r2 : in STD_LOGIC_VECTOR(127 downto 0);
       r3 : in STD_LOGIC_VECTOR(127 downto 0);
       alu_out : out STD_LOGIC_VECTOR(127 downto 0);
       ins_out : out STD_LOGIC_VECTOR(24 downto 0)
  );
end component;
component forwarding_unit
  port (
       ALU_out : in STD_LOGIC_VECTOR(127 downto 0);
       ins : in STD_LOGIC_VECTOR(24 downto 0);
       old_ins : in STD_LOGIC_VECTOR(24 downto 0);
       r1_in : in STD_LOGIC_VECTOR(127 downto 0);
       r2_in : in STD_LOGIC_VECTOR(127 downto 0);
       r3_in : in STD_LOGIC_VECTOR(127 downto 0);
       r1_out : out STD_LOGIC_VECTOR(127 downto 0);
       r2_out : out STD_LOGIC_VECTOR(127 downto 0);
       r3_out : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;
component ins_buffer
  port (
       clk : in STD_LOGIC;
       instructions : in insBuffer;
       ins_out : out STD_LOGIC_VECTOR(24 downto 0)
  );
end component;
component register_file
  port (
       WrData : in STD_LOGIC_VECTOR(127 downto 0);
       clk : in STD_LOGIC;
       ins : in STD_LOGIC_VECTOR(24 downto 0);
       old_ins : in STD_LOGIC_VECTOR(24 downto 0);
       ins_out : out STD_LOGIC_VECTOR(24 downto 0);
       r1 : out STD_LOGIC_VECTOR(127 downto 0);
       r2 : out STD_LOGIC_VECTOR(127 downto 0);
       r3 : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;

----     Constants     -----
constant DANGLING_INPUT_CONSTANT : STD_LOGIC := 'Z';

---- Signal declarations used on the diagram ----

signal NET114 : STD_LOGIC;
signal NET122 : STD_LOGIC;
signal NET134 : STD_LOGIC;
signal NET168 : STD_LOGIC;
signal NET180 : STD_LOGIC;
signal NET210 : STD_LOGIC;
signal NET222 : STD_LOGIC;
signal NET230 : STD_LOGIC;
signal NET238 : STD_LOGIC;
signal NET246 : STD_LOGIC;

---- Declaration for Dangling input ----
signal Dangling_Input_Signal : STD_LOGIC;

---- Declarations for Dangling outputs ----
signal DANGLING_U1_ins_out_23 : STD_LOGIC;
signal DANGLING_U1_ins_out_22 : STD_LOGIC;
signal DANGLING_U1_ins_out_21 : STD_LOGIC;
signal DANGLING_U1_ins_out_20 : STD_LOGIC;
signal DANGLING_U1_ins_out_19 : STD_LOGIC;
signal DANGLING_U1_ins_out_18 : STD_LOGIC;
signal DANGLING_U1_ins_out_17 : STD_LOGIC;
signal DANGLING_U1_ins_out_16 : STD_LOGIC;
signal DANGLING_U1_ins_out_15 : STD_LOGIC;
signal DANGLING_U1_ins_out_14 : STD_LOGIC;
signal DANGLING_U1_ins_out_13 : STD_LOGIC;
signal DANGLING_U1_ins_out_12 : STD_LOGIC;
signal DANGLING_U1_ins_out_11 : STD_LOGIC;
signal DANGLING_U1_ins_out_10 : STD_LOGIC;
signal DANGLING_U1_ins_out_9 : STD_LOGIC;
signal DANGLING_U1_ins_out_8 : STD_LOGIC;
signal DANGLING_U1_ins_out_7 : STD_LOGIC;
signal DANGLING_U1_ins_out_6 : STD_LOGIC;
signal DANGLING_U1_ins_out_5 : STD_LOGIC;
signal DANGLING_U1_ins_out_4 : STD_LOGIC;
signal DANGLING_U1_ins_out_3 : STD_LOGIC;
signal DANGLING_U1_ins_out_2 : STD_LOGIC;
signal DANGLING_U1_ins_out_1 : STD_LOGIC;
signal DANGLING_U1_ins_out_0 : STD_LOGIC;
signal DANGLING_U2_ins_out_23 : STD_LOGIC;
signal DANGLING_U2_ins_out_22 : STD_LOGIC;
signal DANGLING_U2_ins_out_21 : STD_LOGIC;
signal DANGLING_U2_ins_out_20 : STD_LOGIC;
signal DANGLING_U2_ins_out_19 : STD_LOGIC;
signal DANGLING_U2_ins_out_18 : STD_LOGIC;
signal DANGLING_U2_ins_out_17 : STD_LOGIC;
signal DANGLING_U2_ins_out_16 : STD_LOGIC;
signal DANGLING_U2_ins_out_15 : STD_LOGIC;
signal DANGLING_U2_ins_out_14 : STD_LOGIC;
signal DANGLING_U2_ins_out_13 : STD_LOGIC;
signal DANGLING_U2_ins_out_12 : STD_LOGIC;
signal DANGLING_U2_ins_out_11 : STD_LOGIC;
signal DANGLING_U2_ins_out_10 : STD_LOGIC;
signal DANGLING_U2_ins_out_9 : STD_LOGIC;
signal DANGLING_U2_ins_out_8 : STD_LOGIC;
signal DANGLING_U2_ins_out_7 : STD_LOGIC;
signal DANGLING_U2_ins_out_6 : STD_LOGIC;
signal DANGLING_U2_ins_out_5 : STD_LOGIC;
signal DANGLING_U2_ins_out_4 : STD_LOGIC;
signal DANGLING_U2_ins_out_3 : STD_LOGIC;
signal DANGLING_U2_ins_out_2 : STD_LOGIC;
signal DANGLING_U2_ins_out_1 : STD_LOGIC;
signal DANGLING_U2_ins_out_0 : STD_LOGIC;
signal DANGLING_U2_alu_out_126 : STD_LOGIC;
signal DANGLING_U2_alu_out_125 : STD_LOGIC;
signal DANGLING_U2_alu_out_124 : STD_LOGIC;
signal DANGLING_U2_alu_out_123 : STD_LOGIC;
signal DANGLING_U2_alu_out_122 : STD_LOGIC;
signal DANGLING_U2_alu_out_121 : STD_LOGIC;
signal DANGLING_U2_alu_out_120 : STD_LOGIC;
signal DANGLING_U2_alu_out_119 : STD_LOGIC;
signal DANGLING_U2_alu_out_118 : STD_LOGIC;
signal DANGLING_U2_alu_out_117 : STD_LOGIC;
signal DANGLING_U2_alu_out_116 : STD_LOGIC;
signal DANGLING_U2_alu_out_115 : STD_LOGIC;
signal DANGLING_U2_alu_out_114 : STD_LOGIC;
signal DANGLING_U2_alu_out_113 : STD_LOGIC;
signal DANGLING_U2_alu_out_112 : STD_LOGIC;
signal DANGLING_U2_alu_out_111 : STD_LOGIC;
signal DANGLING_U2_alu_out_110 : STD_LOGIC;
signal DANGLING_U2_alu_out_109 : STD_LOGIC;
signal DANGLING_U2_alu_out_108 : STD_LOGIC;
signal DANGLING_U2_alu_out_107 : STD_LOGIC;
signal DANGLING_U2_alu_out_106 : STD_LOGIC;
signal DANGLING_U2_alu_out_105 : STD_LOGIC;
signal DANGLING_U2_alu_out_104 : STD_LOGIC;
signal DANGLING_U2_alu_out_103 : STD_LOGIC;
signal DANGLING_U2_alu_out_102 : STD_LOGIC;
signal DANGLING_U2_alu_out_101 : STD_LOGIC;
signal DANGLING_U2_alu_out_100 : STD_LOGIC;
signal DANGLING_U2_alu_out_99 : STD_LOGIC;
signal DANGLING_U2_alu_out_98 : STD_LOGIC;
signal DANGLING_U2_alu_out_97 : STD_LOGIC;
signal DANGLING_U2_alu_out_96 : STD_LOGIC;
signal DANGLING_U2_alu_out_95 : STD_LOGIC;
signal DANGLING_U2_alu_out_94 : STD_LOGIC;
signal DANGLING_U2_alu_out_93 : STD_LOGIC;
signal DANGLING_U2_alu_out_92 : STD_LOGIC;
signal DANGLING_U2_alu_out_91 : STD_LOGIC;
signal DANGLING_U2_alu_out_90 : STD_LOGIC;
signal DANGLING_U2_alu_out_89 : STD_LOGIC;
signal DANGLING_U2_alu_out_88 : STD_LOGIC;
signal DANGLING_U2_alu_out_87 : STD_LOGIC;
signal DANGLING_U2_alu_out_86 : STD_LOGIC;
signal DANGLING_U2_alu_out_85 : STD_LOGIC;
signal DANGLING_U2_alu_out_84 : STD_LOGIC;
signal DANGLING_U2_alu_out_83 : STD_LOGIC;
signal DANGLING_U2_alu_out_82 : STD_LOGIC;
signal DANGLING_U2_alu_out_81 : STD_LOGIC;
signal DANGLING_U2_alu_out_80 : STD_LOGIC;
signal DANGLING_U2_alu_out_79 : STD_LOGIC;
signal DANGLING_U2_alu_out_78 : STD_LOGIC;
signal DANGLING_U2_alu_out_77 : STD_LOGIC;
signal DANGLING_U2_alu_out_76 : STD_LOGIC;
signal DANGLING_U2_alu_out_75 : STD_LOGIC;
signal DANGLING_U2_alu_out_74 : STD_LOGIC;
signal DANGLING_U2_alu_out_73 : STD_LOGIC;
signal DANGLING_U2_alu_out_72 : STD_LOGIC;
signal DANGLING_U2_alu_out_71 : STD_LOGIC;
signal DANGLING_U2_alu_out_70 : STD_LOGIC;
signal DANGLING_U2_alu_out_69 : STD_LOGIC;
signal DANGLING_U2_alu_out_68 : STD_LOGIC;
signal DANGLING_U2_alu_out_67 : STD_LOGIC;
signal DANGLING_U2_alu_out_66 : STD_LOGIC;
signal DANGLING_U2_alu_out_65 : STD_LOGIC;
signal DANGLING_U2_alu_out_64 : STD_LOGIC;
signal DANGLING_U2_alu_out_63 : STD_LOGIC;
signal DANGLING_U2_alu_out_62 : STD_LOGIC;
signal DANGLING_U2_alu_out_61 : STD_LOGIC;
signal DANGLING_U2_alu_out_60 : STD_LOGIC;
signal DANGLING_U2_alu_out_59 : STD_LOGIC;
signal DANGLING_U2_alu_out_58 : STD_LOGIC;
signal DANGLING_U2_alu_out_57 : STD_LOGIC;
signal DANGLING_U2_alu_out_56 : STD_LOGIC;
signal DANGLING_U2_alu_out_55 : STD_LOGIC;
signal DANGLING_U2_alu_out_54 : STD_LOGIC;
signal DANGLING_U2_alu_out_53 : STD_LOGIC;
signal DANGLING_U2_alu_out_52 : STD_LOGIC;
signal DANGLING_U2_alu_out_51 : STD_LOGIC;
signal DANGLING_U2_alu_out_50 : STD_LOGIC;
signal DANGLING_U2_alu_out_49 : STD_LOGIC;
signal DANGLING_U2_alu_out_48 : STD_LOGIC;
signal DANGLING_U2_alu_out_47 : STD_LOGIC;
signal DANGLING_U2_alu_out_46 : STD_LOGIC;
signal DANGLING_U2_alu_out_45 : STD_LOGIC;
signal DANGLING_U2_alu_out_44 : STD_LOGIC;
signal DANGLING_U2_alu_out_43 : STD_LOGIC;
signal DANGLING_U2_alu_out_42 : STD_LOGIC;
signal DANGLING_U2_alu_out_41 : STD_LOGIC;
signal DANGLING_U2_alu_out_40 : STD_LOGIC;
signal DANGLING_U2_alu_out_39 : STD_LOGIC;
signal DANGLING_U2_alu_out_38 : STD_LOGIC;
signal DANGLING_U2_alu_out_37 : STD_LOGIC;
signal DANGLING_U2_alu_out_36 : STD_LOGIC;
signal DANGLING_U2_alu_out_35 : STD_LOGIC;
signal DANGLING_U2_alu_out_34 : STD_LOGIC;
signal DANGLING_U2_alu_out_33 : STD_LOGIC;
signal DANGLING_U2_alu_out_32 : STD_LOGIC;
signal DANGLING_U2_alu_out_31 : STD_LOGIC;
signal DANGLING_U2_alu_out_30 : STD_LOGIC;
signal DANGLING_U2_alu_out_29 : STD_LOGIC;
signal DANGLING_U2_alu_out_28 : STD_LOGIC;
signal DANGLING_U2_alu_out_27 : STD_LOGIC;
signal DANGLING_U2_alu_out_26 : STD_LOGIC;
signal DANGLING_U2_alu_out_25 : STD_LOGIC;
signal DANGLING_U2_alu_out_24 : STD_LOGIC;
signal DANGLING_U2_alu_out_23 : STD_LOGIC;
signal DANGLING_U2_alu_out_22 : STD_LOGIC;
signal DANGLING_U2_alu_out_21 : STD_LOGIC;
signal DANGLING_U2_alu_out_20 : STD_LOGIC;
signal DANGLING_U2_alu_out_19 : STD_LOGIC;
signal DANGLING_U2_alu_out_18 : STD_LOGIC;
signal DANGLING_U2_alu_out_17 : STD_LOGIC;
signal DANGLING_U2_alu_out_16 : STD_LOGIC;
signal DANGLING_U2_alu_out_15 : STD_LOGIC;
signal DANGLING_U2_alu_out_14 : STD_LOGIC;
signal DANGLING_U2_alu_out_13 : STD_LOGIC;
signal DANGLING_U2_alu_out_12 : STD_LOGIC;
signal DANGLING_U2_alu_out_11 : STD_LOGIC;
signal DANGLING_U2_alu_out_10 : STD_LOGIC;
signal DANGLING_U2_alu_out_9 : STD_LOGIC;
signal DANGLING_U2_alu_out_8 : STD_LOGIC;
signal DANGLING_U2_alu_out_7 : STD_LOGIC;
signal DANGLING_U2_alu_out_6 : STD_LOGIC;
signal DANGLING_U2_alu_out_5 : STD_LOGIC;
signal DANGLING_U2_alu_out_4 : STD_LOGIC;
signal DANGLING_U2_alu_out_3 : STD_LOGIC;
signal DANGLING_U2_alu_out_2 : STD_LOGIC;
signal DANGLING_U2_alu_out_1 : STD_LOGIC;
signal DANGLING_U2_alu_out_0 : STD_LOGIC;
signal DANGLING_U3_r1_out_126 : STD_LOGIC;
signal DANGLING_U3_r1_out_125 : STD_LOGIC;
signal DANGLING_U3_r1_out_124 : STD_LOGIC;
signal DANGLING_U3_r1_out_123 : STD_LOGIC;
signal DANGLING_U3_r1_out_122 : STD_LOGIC;
signal DANGLING_U3_r1_out_121 : STD_LOGIC;
signal DANGLING_U3_r1_out_120 : STD_LOGIC;
signal DANGLING_U3_r1_out_119 : STD_LOGIC;
signal DANGLING_U3_r1_out_118 : STD_LOGIC;
signal DANGLING_U3_r1_out_117 : STD_LOGIC;
signal DANGLING_U3_r1_out_116 : STD_LOGIC;
signal DANGLING_U3_r1_out_115 : STD_LOGIC;
signal DANGLING_U3_r1_out_114 : STD_LOGIC;
signal DANGLING_U3_r1_out_113 : STD_LOGIC;
signal DANGLING_U3_r1_out_112 : STD_LOGIC;
signal DANGLING_U3_r1_out_111 : STD_LOGIC;
signal DANGLING_U3_r1_out_110 : STD_LOGIC;
signal DANGLING_U3_r1_out_109 : STD_LOGIC;
signal DANGLING_U3_r1_out_108 : STD_LOGIC;
signal DANGLING_U3_r1_out_107 : STD_LOGIC;
signal DANGLING_U3_r1_out_106 : STD_LOGIC;
signal DANGLING_U3_r1_out_105 : STD_LOGIC;
signal DANGLING_U3_r1_out_104 : STD_LOGIC;
signal DANGLING_U3_r1_out_103 : STD_LOGIC;
signal DANGLING_U3_r1_out_102 : STD_LOGIC;
signal DANGLING_U3_r1_out_101 : STD_LOGIC;
signal DANGLING_U3_r1_out_100 : STD_LOGIC;
signal DANGLING_U3_r1_out_99 : STD_LOGIC;
signal DANGLING_U3_r1_out_98 : STD_LOGIC;
signal DANGLING_U3_r1_out_97 : STD_LOGIC;
signal DANGLING_U3_r1_out_96 : STD_LOGIC;
signal DANGLING_U3_r1_out_95 : STD_LOGIC;
signal DANGLING_U3_r1_out_94 : STD_LOGIC;
signal DANGLING_U3_r1_out_93 : STD_LOGIC;
signal DANGLING_U3_r1_out_92 : STD_LOGIC;
signal DANGLING_U3_r1_out_91 : STD_LOGIC;
signal DANGLING_U3_r1_out_90 : STD_LOGIC;
signal DANGLING_U3_r1_out_89 : STD_LOGIC;
signal DANGLING_U3_r1_out_88 : STD_LOGIC;
signal DANGLING_U3_r1_out_87 : STD_LOGIC;
signal DANGLING_U3_r1_out_86 : STD_LOGIC;
signal DANGLING_U3_r1_out_85 : STD_LOGIC;
signal DANGLING_U3_r1_out_84 : STD_LOGIC;
signal DANGLING_U3_r1_out_83 : STD_LOGIC;
signal DANGLING_U3_r1_out_82 : STD_LOGIC;
signal DANGLING_U3_r1_out_81 : STD_LOGIC;
signal DANGLING_U3_r1_out_80 : STD_LOGIC;
signal DANGLING_U3_r1_out_79 : STD_LOGIC;
signal DANGLING_U3_r1_out_78 : STD_LOGIC;
signal DANGLING_U3_r1_out_77 : STD_LOGIC;
signal DANGLING_U3_r1_out_76 : STD_LOGIC;
signal DANGLING_U3_r1_out_75 : STD_LOGIC;
signal DANGLING_U3_r1_out_74 : STD_LOGIC;
signal DANGLING_U3_r1_out_73 : STD_LOGIC;
signal DANGLING_U3_r1_out_72 : STD_LOGIC;
signal DANGLING_U3_r1_out_71 : STD_LOGIC;
signal DANGLING_U3_r1_out_70 : STD_LOGIC;
signal DANGLING_U3_r1_out_69 : STD_LOGIC;
signal DANGLING_U3_r1_out_68 : STD_LOGIC;
signal DANGLING_U3_r1_out_67 : STD_LOGIC;
signal DANGLING_U3_r1_out_66 : STD_LOGIC;
signal DANGLING_U3_r1_out_65 : STD_LOGIC;
signal DANGLING_U3_r1_out_64 : STD_LOGIC;
signal DANGLING_U3_r1_out_63 : STD_LOGIC;
signal DANGLING_U3_r1_out_62 : STD_LOGIC;
signal DANGLING_U3_r1_out_61 : STD_LOGIC;
signal DANGLING_U3_r1_out_60 : STD_LOGIC;
signal DANGLING_U3_r1_out_59 : STD_LOGIC;
signal DANGLING_U3_r1_out_58 : STD_LOGIC;
signal DANGLING_U3_r1_out_57 : STD_LOGIC;
signal DANGLING_U3_r1_out_56 : STD_LOGIC;
signal DANGLING_U3_r1_out_55 : STD_LOGIC;
signal DANGLING_U3_r1_out_54 : STD_LOGIC;
signal DANGLING_U3_r1_out_53 : STD_LOGIC;
signal DANGLING_U3_r1_out_52 : STD_LOGIC;
signal DANGLING_U3_r1_out_51 : STD_LOGIC;
signal DANGLING_U3_r1_out_50 : STD_LOGIC;
signal DANGLING_U3_r1_out_49 : STD_LOGIC;
signal DANGLING_U3_r1_out_48 : STD_LOGIC;
signal DANGLING_U3_r1_out_47 : STD_LOGIC;
signal DANGLING_U3_r1_out_46 : STD_LOGIC;
signal DANGLING_U3_r1_out_45 : STD_LOGIC;
signal DANGLING_U3_r1_out_44 : STD_LOGIC;
signal DANGLING_U3_r1_out_43 : STD_LOGIC;
signal DANGLING_U3_r1_out_42 : STD_LOGIC;
signal DANGLING_U3_r1_out_41 : STD_LOGIC;
signal DANGLING_U3_r1_out_40 : STD_LOGIC;
signal DANGLING_U3_r1_out_39 : STD_LOGIC;
signal DANGLING_U3_r1_out_38 : STD_LOGIC;
signal DANGLING_U3_r1_out_37 : STD_LOGIC;
signal DANGLING_U3_r1_out_36 : STD_LOGIC;
signal DANGLING_U3_r1_out_35 : STD_LOGIC;
signal DANGLING_U3_r1_out_34 : STD_LOGIC;
signal DANGLING_U3_r1_out_33 : STD_LOGIC;
signal DANGLING_U3_r1_out_32 : STD_LOGIC;
signal DANGLING_U3_r1_out_31 : STD_LOGIC;
signal DANGLING_U3_r1_out_30 : STD_LOGIC;
signal DANGLING_U3_r1_out_29 : STD_LOGIC;
signal DANGLING_U3_r1_out_28 : STD_LOGIC;
signal DANGLING_U3_r1_out_27 : STD_LOGIC;
signal DANGLING_U3_r1_out_26 : STD_LOGIC;
signal DANGLING_U3_r1_out_25 : STD_LOGIC;
signal DANGLING_U3_r1_out_24 : STD_LOGIC;
signal DANGLING_U3_r1_out_23 : STD_LOGIC;
signal DANGLING_U3_r1_out_22 : STD_LOGIC;
signal DANGLING_U3_r1_out_21 : STD_LOGIC;
signal DANGLING_U3_r1_out_20 : STD_LOGIC;
signal DANGLING_U3_r1_out_19 : STD_LOGIC;
signal DANGLING_U3_r1_out_18 : STD_LOGIC;
signal DANGLING_U3_r1_out_17 : STD_LOGIC;
signal DANGLING_U3_r1_out_16 : STD_LOGIC;
signal DANGLING_U3_r1_out_15 : STD_LOGIC;
signal DANGLING_U3_r1_out_14 : STD_LOGIC;
signal DANGLING_U3_r1_out_13 : STD_LOGIC;
signal DANGLING_U3_r1_out_12 : STD_LOGIC;
signal DANGLING_U3_r1_out_11 : STD_LOGIC;
signal DANGLING_U3_r1_out_10 : STD_LOGIC;
signal DANGLING_U3_r1_out_9 : STD_LOGIC;
signal DANGLING_U3_r1_out_8 : STD_LOGIC;
signal DANGLING_U3_r1_out_7 : STD_LOGIC;
signal DANGLING_U3_r1_out_6 : STD_LOGIC;
signal DANGLING_U3_r1_out_5 : STD_LOGIC;
signal DANGLING_U3_r1_out_4 : STD_LOGIC;
signal DANGLING_U3_r1_out_3 : STD_LOGIC;
signal DANGLING_U3_r1_out_2 : STD_LOGIC;
signal DANGLING_U3_r1_out_1 : STD_LOGIC;
signal DANGLING_U3_r1_out_0 : STD_LOGIC;
signal DANGLING_U3_r2_out_126 : STD_LOGIC;
signal DANGLING_U3_r2_out_125 : STD_LOGIC;
signal DANGLING_U3_r2_out_124 : STD_LOGIC;
signal DANGLING_U3_r2_out_123 : STD_LOGIC;
signal DANGLING_U3_r2_out_122 : STD_LOGIC;
signal DANGLING_U3_r2_out_121 : STD_LOGIC;
signal DANGLING_U3_r2_out_120 : STD_LOGIC;
signal DANGLING_U3_r2_out_119 : STD_LOGIC;
signal DANGLING_U3_r2_out_118 : STD_LOGIC;
signal DANGLING_U3_r2_out_117 : STD_LOGIC;
signal DANGLING_U3_r2_out_116 : STD_LOGIC;
signal DANGLING_U3_r2_out_115 : STD_LOGIC;
signal DANGLING_U3_r2_out_114 : STD_LOGIC;
signal DANGLING_U3_r2_out_113 : STD_LOGIC;
signal DANGLING_U3_r2_out_112 : STD_LOGIC;
signal DANGLING_U3_r2_out_111 : STD_LOGIC;
signal DANGLING_U3_r2_out_110 : STD_LOGIC;
signal DANGLING_U3_r2_out_109 : STD_LOGIC;
signal DANGLING_U3_r2_out_108 : STD_LOGIC;
signal DANGLING_U3_r2_out_107 : STD_LOGIC;
signal DANGLING_U3_r2_out_106 : STD_LOGIC;
signal DANGLING_U3_r2_out_105 : STD_LOGIC;
signal DANGLING_U3_r2_out_104 : STD_LOGIC;
signal DANGLING_U3_r2_out_103 : STD_LOGIC;
signal DANGLING_U3_r2_out_102 : STD_LOGIC;
signal DANGLING_U3_r2_out_101 : STD_LOGIC;
signal DANGLING_U3_r2_out_100 : STD_LOGIC;
signal DANGLING_U3_r2_out_99 : STD_LOGIC;
signal DANGLING_U3_r2_out_98 : STD_LOGIC;
signal DANGLING_U3_r2_out_97 : STD_LOGIC;
signal DANGLING_U3_r2_out_96 : STD_LOGIC;
signal DANGLING_U3_r2_out_95 : STD_LOGIC;
signal DANGLING_U3_r2_out_94 : STD_LOGIC;
signal DANGLING_U3_r2_out_93 : STD_LOGIC;
signal DANGLING_U3_r2_out_92 : STD_LOGIC;
signal DANGLING_U3_r2_out_91 : STD_LOGIC;
signal DANGLING_U3_r2_out_90 : STD_LOGIC;
signal DANGLING_U3_r2_out_89 : STD_LOGIC;
signal DANGLING_U3_r2_out_88 : STD_LOGIC;
signal DANGLING_U3_r2_out_87 : STD_LOGIC;
signal DANGLING_U3_r2_out_86 : STD_LOGIC;
signal DANGLING_U3_r2_out_85 : STD_LOGIC;
signal DANGLING_U3_r2_out_84 : STD_LOGIC;
signal DANGLING_U3_r2_out_83 : STD_LOGIC;
signal DANGLING_U3_r2_out_82 : STD_LOGIC;
signal DANGLING_U3_r2_out_81 : STD_LOGIC;
signal DANGLING_U3_r2_out_80 : STD_LOGIC;
signal DANGLING_U3_r2_out_79 : STD_LOGIC;
signal DANGLING_U3_r2_out_78 : STD_LOGIC;
signal DANGLING_U3_r2_out_77 : STD_LOGIC;
signal DANGLING_U3_r2_out_76 : STD_LOGIC;
signal DANGLING_U3_r2_out_75 : STD_LOGIC;
signal DANGLING_U3_r2_out_74 : STD_LOGIC;
signal DANGLING_U3_r2_out_73 : STD_LOGIC;
signal DANGLING_U3_r2_out_72 : STD_LOGIC;
signal DANGLING_U3_r2_out_71 : STD_LOGIC;
signal DANGLING_U3_r2_out_70 : STD_LOGIC;
signal DANGLING_U3_r2_out_69 : STD_LOGIC;
signal DANGLING_U3_r2_out_68 : STD_LOGIC;
signal DANGLING_U3_r2_out_67 : STD_LOGIC;
signal DANGLING_U3_r2_out_66 : STD_LOGIC;
signal DANGLING_U3_r2_out_65 : STD_LOGIC;
signal DANGLING_U3_r2_out_64 : STD_LOGIC;
signal DANGLING_U3_r2_out_63 : STD_LOGIC;
signal DANGLING_U3_r2_out_62 : STD_LOGIC;
signal DANGLING_U3_r2_out_61 : STD_LOGIC;
signal DANGLING_U3_r2_out_60 : STD_LOGIC;
signal DANGLING_U3_r2_out_59 : STD_LOGIC;
signal DANGLING_U3_r2_out_58 : STD_LOGIC;
signal DANGLING_U3_r2_out_57 : STD_LOGIC;
signal DANGLING_U3_r2_out_56 : STD_LOGIC;
signal DANGLING_U3_r2_out_55 : STD_LOGIC;
signal DANGLING_U3_r2_out_54 : STD_LOGIC;
signal DANGLING_U3_r2_out_53 : STD_LOGIC;
signal DANGLING_U3_r2_out_52 : STD_LOGIC;
signal DANGLING_U3_r2_out_51 : STD_LOGIC;
signal DANGLING_U3_r2_out_50 : STD_LOGIC;
signal DANGLING_U3_r2_out_49 : STD_LOGIC;
signal DANGLING_U3_r2_out_48 : STD_LOGIC;
signal DANGLING_U3_r2_out_47 : STD_LOGIC;
signal DANGLING_U3_r2_out_46 : STD_LOGIC;
signal DANGLING_U3_r2_out_45 : STD_LOGIC;
signal DANGLING_U3_r2_out_44 : STD_LOGIC;
signal DANGLING_U3_r2_out_43 : STD_LOGIC;
signal DANGLING_U3_r2_out_42 : STD_LOGIC;
signal DANGLING_U3_r2_out_41 : STD_LOGIC;
signal DANGLING_U3_r2_out_40 : STD_LOGIC;
signal DANGLING_U3_r2_out_39 : STD_LOGIC;
signal DANGLING_U3_r2_out_38 : STD_LOGIC;
signal DANGLING_U3_r2_out_37 : STD_LOGIC;
signal DANGLING_U3_r2_out_36 : STD_LOGIC;
signal DANGLING_U3_r2_out_35 : STD_LOGIC;
signal DANGLING_U3_r2_out_34 : STD_LOGIC;
signal DANGLING_U3_r2_out_33 : STD_LOGIC;
signal DANGLING_U3_r2_out_32 : STD_LOGIC;
signal DANGLING_U3_r2_out_31 : STD_LOGIC;
signal DANGLING_U3_r2_out_30 : STD_LOGIC;
signal DANGLING_U3_r2_out_29 : STD_LOGIC;
signal DANGLING_U3_r2_out_28 : STD_LOGIC;
signal DANGLING_U3_r2_out_27 : STD_LOGIC;
signal DANGLING_U3_r2_out_26 : STD_LOGIC;
signal DANGLING_U3_r2_out_25 : STD_LOGIC;
signal DANGLING_U3_r2_out_24 : STD_LOGIC;
signal DANGLING_U3_r2_out_23 : STD_LOGIC;
signal DANGLING_U3_r2_out_22 : STD_LOGIC;
signal DANGLING_U3_r2_out_21 : STD_LOGIC;
signal DANGLING_U3_r2_out_20 : STD_LOGIC;
signal DANGLING_U3_r2_out_19 : STD_LOGIC;
signal DANGLING_U3_r2_out_18 : STD_LOGIC;
signal DANGLING_U3_r2_out_17 : STD_LOGIC;
signal DANGLING_U3_r2_out_16 : STD_LOGIC;
signal DANGLING_U3_r2_out_15 : STD_LOGIC;
signal DANGLING_U3_r2_out_14 : STD_LOGIC;
signal DANGLING_U3_r2_out_13 : STD_LOGIC;
signal DANGLING_U3_r2_out_12 : STD_LOGIC;
signal DANGLING_U3_r2_out_11 : STD_LOGIC;
signal DANGLING_U3_r2_out_10 : STD_LOGIC;
signal DANGLING_U3_r2_out_9 : STD_LOGIC;
signal DANGLING_U3_r2_out_8 : STD_LOGIC;
signal DANGLING_U3_r2_out_7 : STD_LOGIC;
signal DANGLING_U3_r2_out_6 : STD_LOGIC;
signal DANGLING_U3_r2_out_5 : STD_LOGIC;
signal DANGLING_U3_r2_out_4 : STD_LOGIC;
signal DANGLING_U3_r2_out_3 : STD_LOGIC;
signal DANGLING_U3_r2_out_2 : STD_LOGIC;
signal DANGLING_U3_r2_out_1 : STD_LOGIC;
signal DANGLING_U3_r2_out_0 : STD_LOGIC;
signal DANGLING_U3_r3_out_126 : STD_LOGIC;
signal DANGLING_U3_r3_out_125 : STD_LOGIC;
signal DANGLING_U3_r3_out_124 : STD_LOGIC;
signal DANGLING_U3_r3_out_123 : STD_LOGIC;
signal DANGLING_U3_r3_out_122 : STD_LOGIC;
signal DANGLING_U3_r3_out_121 : STD_LOGIC;
signal DANGLING_U3_r3_out_120 : STD_LOGIC;
signal DANGLING_U3_r3_out_119 : STD_LOGIC;
signal DANGLING_U3_r3_out_118 : STD_LOGIC;
signal DANGLING_U3_r3_out_117 : STD_LOGIC;
signal DANGLING_U3_r3_out_116 : STD_LOGIC;
signal DANGLING_U3_r3_out_115 : STD_LOGIC;
signal DANGLING_U3_r3_out_114 : STD_LOGIC;
signal DANGLING_U3_r3_out_113 : STD_LOGIC;
signal DANGLING_U3_r3_out_112 : STD_LOGIC;
signal DANGLING_U3_r3_out_111 : STD_LOGIC;
signal DANGLING_U3_r3_out_110 : STD_LOGIC;
signal DANGLING_U3_r3_out_109 : STD_LOGIC;
signal DANGLING_U3_r3_out_108 : STD_LOGIC;
signal DANGLING_U3_r3_out_107 : STD_LOGIC;
signal DANGLING_U3_r3_out_106 : STD_LOGIC;
signal DANGLING_U3_r3_out_105 : STD_LOGIC;
signal DANGLING_U3_r3_out_104 : STD_LOGIC;
signal DANGLING_U3_r3_out_103 : STD_LOGIC;
signal DANGLING_U3_r3_out_102 : STD_LOGIC;
signal DANGLING_U3_r3_out_101 : STD_LOGIC;
signal DANGLING_U3_r3_out_100 : STD_LOGIC;
signal DANGLING_U3_r3_out_99 : STD_LOGIC;
signal DANGLING_U3_r3_out_98 : STD_LOGIC;
signal DANGLING_U3_r3_out_97 : STD_LOGIC;
signal DANGLING_U3_r3_out_96 : STD_LOGIC;
signal DANGLING_U3_r3_out_95 : STD_LOGIC;
signal DANGLING_U3_r3_out_94 : STD_LOGIC;
signal DANGLING_U3_r3_out_93 : STD_LOGIC;
signal DANGLING_U3_r3_out_92 : STD_LOGIC;
signal DANGLING_U3_r3_out_91 : STD_LOGIC;
signal DANGLING_U3_r3_out_90 : STD_LOGIC;
signal DANGLING_U3_r3_out_89 : STD_LOGIC;
signal DANGLING_U3_r3_out_88 : STD_LOGIC;
signal DANGLING_U3_r3_out_87 : STD_LOGIC;
signal DANGLING_U3_r3_out_86 : STD_LOGIC;
signal DANGLING_U3_r3_out_85 : STD_LOGIC;
signal DANGLING_U3_r3_out_84 : STD_LOGIC;
signal DANGLING_U3_r3_out_83 : STD_LOGIC;
signal DANGLING_U3_r3_out_82 : STD_LOGIC;
signal DANGLING_U3_r3_out_81 : STD_LOGIC;
signal DANGLING_U3_r3_out_80 : STD_LOGIC;
signal DANGLING_U3_r3_out_79 : STD_LOGIC;
signal DANGLING_U3_r3_out_78 : STD_LOGIC;
signal DANGLING_U3_r3_out_77 : STD_LOGIC;
signal DANGLING_U3_r3_out_76 : STD_LOGIC;
signal DANGLING_U3_r3_out_75 : STD_LOGIC;
signal DANGLING_U3_r3_out_74 : STD_LOGIC;
signal DANGLING_U3_r3_out_73 : STD_LOGIC;
signal DANGLING_U3_r3_out_72 : STD_LOGIC;
signal DANGLING_U3_r3_out_71 : STD_LOGIC;
signal DANGLING_U3_r3_out_70 : STD_LOGIC;
signal DANGLING_U3_r3_out_69 : STD_LOGIC;
signal DANGLING_U3_r3_out_68 : STD_LOGIC;
signal DANGLING_U3_r3_out_67 : STD_LOGIC;
signal DANGLING_U3_r3_out_66 : STD_LOGIC;
signal DANGLING_U3_r3_out_65 : STD_LOGIC;
signal DANGLING_U3_r3_out_64 : STD_LOGIC;
signal DANGLING_U3_r3_out_63 : STD_LOGIC;
signal DANGLING_U3_r3_out_62 : STD_LOGIC;
signal DANGLING_U3_r3_out_61 : STD_LOGIC;
signal DANGLING_U3_r3_out_60 : STD_LOGIC;
signal DANGLING_U3_r3_out_59 : STD_LOGIC;
signal DANGLING_U3_r3_out_58 : STD_LOGIC;
signal DANGLING_U3_r3_out_57 : STD_LOGIC;
signal DANGLING_U3_r3_out_56 : STD_LOGIC;
signal DANGLING_U3_r3_out_55 : STD_LOGIC;
signal DANGLING_U3_r3_out_54 : STD_LOGIC;
signal DANGLING_U3_r3_out_53 : STD_LOGIC;
signal DANGLING_U3_r3_out_52 : STD_LOGIC;
signal DANGLING_U3_r3_out_51 : STD_LOGIC;
signal DANGLING_U3_r3_out_50 : STD_LOGIC;
signal DANGLING_U3_r3_out_49 : STD_LOGIC;
signal DANGLING_U3_r3_out_48 : STD_LOGIC;
signal DANGLING_U3_r3_out_47 : STD_LOGIC;
signal DANGLING_U3_r3_out_46 : STD_LOGIC;
signal DANGLING_U3_r3_out_45 : STD_LOGIC;
signal DANGLING_U3_r3_out_44 : STD_LOGIC;
signal DANGLING_U3_r3_out_43 : STD_LOGIC;
signal DANGLING_U3_r3_out_42 : STD_LOGIC;
signal DANGLING_U3_r3_out_41 : STD_LOGIC;
signal DANGLING_U3_r3_out_40 : STD_LOGIC;
signal DANGLING_U3_r3_out_39 : STD_LOGIC;
signal DANGLING_U3_r3_out_38 : STD_LOGIC;
signal DANGLING_U3_r3_out_37 : STD_LOGIC;
signal DANGLING_U3_r3_out_36 : STD_LOGIC;
signal DANGLING_U3_r3_out_35 : STD_LOGIC;
signal DANGLING_U3_r3_out_34 : STD_LOGIC;
signal DANGLING_U3_r3_out_33 : STD_LOGIC;
signal DANGLING_U3_r3_out_32 : STD_LOGIC;
signal DANGLING_U3_r3_out_31 : STD_LOGIC;
signal DANGLING_U3_r3_out_30 : STD_LOGIC;
signal DANGLING_U3_r3_out_29 : STD_LOGIC;
signal DANGLING_U3_r3_out_28 : STD_LOGIC;
signal DANGLING_U3_r3_out_27 : STD_LOGIC;
signal DANGLING_U3_r3_out_26 : STD_LOGIC;
signal DANGLING_U3_r3_out_25 : STD_LOGIC;
signal DANGLING_U3_r3_out_24 : STD_LOGIC;
signal DANGLING_U3_r3_out_23 : STD_LOGIC;
signal DANGLING_U3_r3_out_22 : STD_LOGIC;
signal DANGLING_U3_r3_out_21 : STD_LOGIC;
signal DANGLING_U3_r3_out_20 : STD_LOGIC;
signal DANGLING_U3_r3_out_19 : STD_LOGIC;
signal DANGLING_U3_r3_out_18 : STD_LOGIC;
signal DANGLING_U3_r3_out_17 : STD_LOGIC;
signal DANGLING_U3_r3_out_16 : STD_LOGIC;
signal DANGLING_U3_r3_out_15 : STD_LOGIC;
signal DANGLING_U3_r3_out_14 : STD_LOGIC;
signal DANGLING_U3_r3_out_13 : STD_LOGIC;
signal DANGLING_U3_r3_out_12 : STD_LOGIC;
signal DANGLING_U3_r3_out_11 : STD_LOGIC;
signal DANGLING_U3_r3_out_10 : STD_LOGIC;
signal DANGLING_U3_r3_out_9 : STD_LOGIC;
signal DANGLING_U3_r3_out_8 : STD_LOGIC;
signal DANGLING_U3_r3_out_7 : STD_LOGIC;
signal DANGLING_U3_r3_out_6 : STD_LOGIC;
signal DANGLING_U3_r3_out_5 : STD_LOGIC;
signal DANGLING_U3_r3_out_4 : STD_LOGIC;
signal DANGLING_U3_r3_out_3 : STD_LOGIC;
signal DANGLING_U3_r3_out_2 : STD_LOGIC;
signal DANGLING_U3_r3_out_1 : STD_LOGIC;
signal DANGLING_U3_r3_out_0 : STD_LOGIC;
signal DANGLING_U5_r1_126 : STD_LOGIC;
signal DANGLING_U5_r1_125 : STD_LOGIC;
signal DANGLING_U5_r1_124 : STD_LOGIC;
signal DANGLING_U5_r1_123 : STD_LOGIC;
signal DANGLING_U5_r1_122 : STD_LOGIC;
signal DANGLING_U5_r1_121 : STD_LOGIC;
signal DANGLING_U5_r1_120 : STD_LOGIC;
signal DANGLING_U5_r1_119 : STD_LOGIC;
signal DANGLING_U5_r1_118 : STD_LOGIC;
signal DANGLING_U5_r1_117 : STD_LOGIC;
signal DANGLING_U5_r1_116 : STD_LOGIC;
signal DANGLING_U5_r1_115 : STD_LOGIC;
signal DANGLING_U5_r1_114 : STD_LOGIC;
signal DANGLING_U5_r1_113 : STD_LOGIC;
signal DANGLING_U5_r1_112 : STD_LOGIC;
signal DANGLING_U5_r1_111 : STD_LOGIC;
signal DANGLING_U5_r1_110 : STD_LOGIC;
signal DANGLING_U5_r1_109 : STD_LOGIC;
signal DANGLING_U5_r1_108 : STD_LOGIC;
signal DANGLING_U5_r1_107 : STD_LOGIC;
signal DANGLING_U5_r1_106 : STD_LOGIC;
signal DANGLING_U5_r1_105 : STD_LOGIC;
signal DANGLING_U5_r1_104 : STD_LOGIC;
signal DANGLING_U5_r1_103 : STD_LOGIC;
signal DANGLING_U5_r1_102 : STD_LOGIC;
signal DANGLING_U5_r1_101 : STD_LOGIC;
signal DANGLING_U5_r1_100 : STD_LOGIC;
signal DANGLING_U5_r1_99 : STD_LOGIC;
signal DANGLING_U5_r1_98 : STD_LOGIC;
signal DANGLING_U5_r1_97 : STD_LOGIC;
signal DANGLING_U5_r1_96 : STD_LOGIC;
signal DANGLING_U5_r1_95 : STD_LOGIC;
signal DANGLING_U5_r1_94 : STD_LOGIC;
signal DANGLING_U5_r1_93 : STD_LOGIC;
signal DANGLING_U5_r1_92 : STD_LOGIC;
signal DANGLING_U5_r1_91 : STD_LOGIC;
signal DANGLING_U5_r1_90 : STD_LOGIC;
signal DANGLING_U5_r1_89 : STD_LOGIC;
signal DANGLING_U5_r1_88 : STD_LOGIC;
signal DANGLING_U5_r1_87 : STD_LOGIC;
signal DANGLING_U5_r1_86 : STD_LOGIC;
signal DANGLING_U5_r1_85 : STD_LOGIC;
signal DANGLING_U5_r1_84 : STD_LOGIC;
signal DANGLING_U5_r1_83 : STD_LOGIC;
signal DANGLING_U5_r1_82 : STD_LOGIC;
signal DANGLING_U5_r1_81 : STD_LOGIC;
signal DANGLING_U5_r1_80 : STD_LOGIC;
signal DANGLING_U5_r1_79 : STD_LOGIC;
signal DANGLING_U5_r1_78 : STD_LOGIC;
signal DANGLING_U5_r1_77 : STD_LOGIC;
signal DANGLING_U5_r1_76 : STD_LOGIC;
signal DANGLING_U5_r1_75 : STD_LOGIC;
signal DANGLING_U5_r1_74 : STD_LOGIC;
signal DANGLING_U5_r1_73 : STD_LOGIC;
signal DANGLING_U5_r1_72 : STD_LOGIC;
signal DANGLING_U5_r1_71 : STD_LOGIC;
signal DANGLING_U5_r1_70 : STD_LOGIC;
signal DANGLING_U5_r1_69 : STD_LOGIC;
signal DANGLING_U5_r1_68 : STD_LOGIC;
signal DANGLING_U5_r1_67 : STD_LOGIC;
signal DANGLING_U5_r1_66 : STD_LOGIC;
signal DANGLING_U5_r1_65 : STD_LOGIC;
signal DANGLING_U5_r1_64 : STD_LOGIC;
signal DANGLING_U5_r1_63 : STD_LOGIC;
signal DANGLING_U5_r1_62 : STD_LOGIC;
signal DANGLING_U5_r1_61 : STD_LOGIC;
signal DANGLING_U5_r1_60 : STD_LOGIC;
signal DANGLING_U5_r1_59 : STD_LOGIC;
signal DANGLING_U5_r1_58 : STD_LOGIC;
signal DANGLING_U5_r1_57 : STD_LOGIC;
signal DANGLING_U5_r1_56 : STD_LOGIC;
signal DANGLING_U5_r1_55 : STD_LOGIC;
signal DANGLING_U5_r1_54 : STD_LOGIC;
signal DANGLING_U5_r1_53 : STD_LOGIC;
signal DANGLING_U5_r1_52 : STD_LOGIC;
signal DANGLING_U5_r1_51 : STD_LOGIC;
signal DANGLING_U5_r1_50 : STD_LOGIC;
signal DANGLING_U5_r1_49 : STD_LOGIC;
signal DANGLING_U5_r1_48 : STD_LOGIC;
signal DANGLING_U5_r1_47 : STD_LOGIC;
signal DANGLING_U5_r1_46 : STD_LOGIC;
signal DANGLING_U5_r1_45 : STD_LOGIC;
signal DANGLING_U5_r1_44 : STD_LOGIC;
signal DANGLING_U5_r1_43 : STD_LOGIC;
signal DANGLING_U5_r1_42 : STD_LOGIC;
signal DANGLING_U5_r1_41 : STD_LOGIC;
signal DANGLING_U5_r1_40 : STD_LOGIC;
signal DANGLING_U5_r1_39 : STD_LOGIC;
signal DANGLING_U5_r1_38 : STD_LOGIC;
signal DANGLING_U5_r1_37 : STD_LOGIC;
signal DANGLING_U5_r1_36 : STD_LOGIC;
signal DANGLING_U5_r1_35 : STD_LOGIC;
signal DANGLING_U5_r1_34 : STD_LOGIC;
signal DANGLING_U5_r1_33 : STD_LOGIC;
signal DANGLING_U5_r1_32 : STD_LOGIC;
signal DANGLING_U5_r1_31 : STD_LOGIC;
signal DANGLING_U5_r1_30 : STD_LOGIC;
signal DANGLING_U5_r1_29 : STD_LOGIC;
signal DANGLING_U5_r1_28 : STD_LOGIC;
signal DANGLING_U5_r1_27 : STD_LOGIC;
signal DANGLING_U5_r1_26 : STD_LOGIC;
signal DANGLING_U5_r1_25 : STD_LOGIC;
signal DANGLING_U5_r1_24 : STD_LOGIC;
signal DANGLING_U5_r1_23 : STD_LOGIC;
signal DANGLING_U5_r1_22 : STD_LOGIC;
signal DANGLING_U5_r1_21 : STD_LOGIC;
signal DANGLING_U5_r1_20 : STD_LOGIC;
signal DANGLING_U5_r1_19 : STD_LOGIC;
signal DANGLING_U5_r1_18 : STD_LOGIC;
signal DANGLING_U5_r1_17 : STD_LOGIC;
signal DANGLING_U5_r1_16 : STD_LOGIC;
signal DANGLING_U5_r1_15 : STD_LOGIC;
signal DANGLING_U5_r1_14 : STD_LOGIC;
signal DANGLING_U5_r1_13 : STD_LOGIC;
signal DANGLING_U5_r1_12 : STD_LOGIC;
signal DANGLING_U5_r1_11 : STD_LOGIC;
signal DANGLING_U5_r1_10 : STD_LOGIC;
signal DANGLING_U5_r1_9 : STD_LOGIC;
signal DANGLING_U5_r1_8 : STD_LOGIC;
signal DANGLING_U5_r1_7 : STD_LOGIC;
signal DANGLING_U5_r1_6 : STD_LOGIC;
signal DANGLING_U5_r1_5 : STD_LOGIC;
signal DANGLING_U5_r1_4 : STD_LOGIC;
signal DANGLING_U5_r1_3 : STD_LOGIC;
signal DANGLING_U5_r1_2 : STD_LOGIC;
signal DANGLING_U5_r1_1 : STD_LOGIC;
signal DANGLING_U5_r1_0 : STD_LOGIC;
signal DANGLING_U5_r2_126 : STD_LOGIC;
signal DANGLING_U5_r2_125 : STD_LOGIC;
signal DANGLING_U5_r2_124 : STD_LOGIC;
signal DANGLING_U5_r2_123 : STD_LOGIC;
signal DANGLING_U5_r2_122 : STD_LOGIC;
signal DANGLING_U5_r2_121 : STD_LOGIC;
signal DANGLING_U5_r2_120 : STD_LOGIC;
signal DANGLING_U5_r2_119 : STD_LOGIC;
signal DANGLING_U5_r2_118 : STD_LOGIC;
signal DANGLING_U5_r2_117 : STD_LOGIC;
signal DANGLING_U5_r2_116 : STD_LOGIC;
signal DANGLING_U5_r2_115 : STD_LOGIC;
signal DANGLING_U5_r2_114 : STD_LOGIC;
signal DANGLING_U5_r2_113 : STD_LOGIC;
signal DANGLING_U5_r2_112 : STD_LOGIC;
signal DANGLING_U5_r2_111 : STD_LOGIC;
signal DANGLING_U5_r2_110 : STD_LOGIC;
signal DANGLING_U5_r2_109 : STD_LOGIC;
signal DANGLING_U5_r2_108 : STD_LOGIC;
signal DANGLING_U5_r2_107 : STD_LOGIC;
signal DANGLING_U5_r2_106 : STD_LOGIC;
signal DANGLING_U5_r2_105 : STD_LOGIC;
signal DANGLING_U5_r2_104 : STD_LOGIC;
signal DANGLING_U5_r2_103 : STD_LOGIC;
signal DANGLING_U5_r2_102 : STD_LOGIC;
signal DANGLING_U5_r2_101 : STD_LOGIC;
signal DANGLING_U5_r2_100 : STD_LOGIC;
signal DANGLING_U5_r2_99 : STD_LOGIC;
signal DANGLING_U5_r2_98 : STD_LOGIC;
signal DANGLING_U5_r2_97 : STD_LOGIC;
signal DANGLING_U5_r2_96 : STD_LOGIC;
signal DANGLING_U5_r2_95 : STD_LOGIC;
signal DANGLING_U5_r2_94 : STD_LOGIC;
signal DANGLING_U5_r2_93 : STD_LOGIC;
signal DANGLING_U5_r2_92 : STD_LOGIC;
signal DANGLING_U5_r2_91 : STD_LOGIC;
signal DANGLING_U5_r2_90 : STD_LOGIC;
signal DANGLING_U5_r2_89 : STD_LOGIC;
signal DANGLING_U5_r2_88 : STD_LOGIC;
signal DANGLING_U5_r2_87 : STD_LOGIC;
signal DANGLING_U5_r2_86 : STD_LOGIC;
signal DANGLING_U5_r2_85 : STD_LOGIC;
signal DANGLING_U5_r2_84 : STD_LOGIC;
signal DANGLING_U5_r2_83 : STD_LOGIC;
signal DANGLING_U5_r2_82 : STD_LOGIC;
signal DANGLING_U5_r2_81 : STD_LOGIC;
signal DANGLING_U5_r2_80 : STD_LOGIC;
signal DANGLING_U5_r2_79 : STD_LOGIC;
signal DANGLING_U5_r2_78 : STD_LOGIC;
signal DANGLING_U5_r2_77 : STD_LOGIC;
signal DANGLING_U5_r2_76 : STD_LOGIC;
signal DANGLING_U5_r2_75 : STD_LOGIC;
signal DANGLING_U5_r2_74 : STD_LOGIC;
signal DANGLING_U5_r2_73 : STD_LOGIC;
signal DANGLING_U5_r2_72 : STD_LOGIC;
signal DANGLING_U5_r2_71 : STD_LOGIC;
signal DANGLING_U5_r2_70 : STD_LOGIC;
signal DANGLING_U5_r2_69 : STD_LOGIC;
signal DANGLING_U5_r2_68 : STD_LOGIC;
signal DANGLING_U5_r2_67 : STD_LOGIC;
signal DANGLING_U5_r2_66 : STD_LOGIC;
signal DANGLING_U5_r2_65 : STD_LOGIC;
signal DANGLING_U5_r2_64 : STD_LOGIC;
signal DANGLING_U5_r2_63 : STD_LOGIC;
signal DANGLING_U5_r2_62 : STD_LOGIC;
signal DANGLING_U5_r2_61 : STD_LOGIC;
signal DANGLING_U5_r2_60 : STD_LOGIC;
signal DANGLING_U5_r2_59 : STD_LOGIC;
signal DANGLING_U5_r2_58 : STD_LOGIC;
signal DANGLING_U5_r2_57 : STD_LOGIC;
signal DANGLING_U5_r2_56 : STD_LOGIC;
signal DANGLING_U5_r2_55 : STD_LOGIC;
signal DANGLING_U5_r2_54 : STD_LOGIC;
signal DANGLING_U5_r2_53 : STD_LOGIC;
signal DANGLING_U5_r2_52 : STD_LOGIC;
signal DANGLING_U5_r2_51 : STD_LOGIC;
signal DANGLING_U5_r2_50 : STD_LOGIC;
signal DANGLING_U5_r2_49 : STD_LOGIC;
signal DANGLING_U5_r2_48 : STD_LOGIC;
signal DANGLING_U5_r2_47 : STD_LOGIC;
signal DANGLING_U5_r2_46 : STD_LOGIC;
signal DANGLING_U5_r2_45 : STD_LOGIC;
signal DANGLING_U5_r2_44 : STD_LOGIC;
signal DANGLING_U5_r2_43 : STD_LOGIC;
signal DANGLING_U5_r2_42 : STD_LOGIC;
signal DANGLING_U5_r2_41 : STD_LOGIC;
signal DANGLING_U5_r2_40 : STD_LOGIC;
signal DANGLING_U5_r2_39 : STD_LOGIC;
signal DANGLING_U5_r2_38 : STD_LOGIC;
signal DANGLING_U5_r2_37 : STD_LOGIC;
signal DANGLING_U5_r2_36 : STD_LOGIC;
signal DANGLING_U5_r2_35 : STD_LOGIC;
signal DANGLING_U5_r2_34 : STD_LOGIC;
signal DANGLING_U5_r2_33 : STD_LOGIC;
signal DANGLING_U5_r2_32 : STD_LOGIC;
signal DANGLING_U5_r2_31 : STD_LOGIC;
signal DANGLING_U5_r2_30 : STD_LOGIC;
signal DANGLING_U5_r2_29 : STD_LOGIC;
signal DANGLING_U5_r2_28 : STD_LOGIC;
signal DANGLING_U5_r2_27 : STD_LOGIC;
signal DANGLING_U5_r2_26 : STD_LOGIC;
signal DANGLING_U5_r2_25 : STD_LOGIC;
signal DANGLING_U5_r2_24 : STD_LOGIC;
signal DANGLING_U5_r2_23 : STD_LOGIC;
signal DANGLING_U5_r2_22 : STD_LOGIC;
signal DANGLING_U5_r2_21 : STD_LOGIC;
signal DANGLING_U5_r2_20 : STD_LOGIC;
signal DANGLING_U5_r2_19 : STD_LOGIC;
signal DANGLING_U5_r2_18 : STD_LOGIC;
signal DANGLING_U5_r2_17 : STD_LOGIC;
signal DANGLING_U5_r2_16 : STD_LOGIC;
signal DANGLING_U5_r2_15 : STD_LOGIC;
signal DANGLING_U5_r2_14 : STD_LOGIC;
signal DANGLING_U5_r2_13 : STD_LOGIC;
signal DANGLING_U5_r2_12 : STD_LOGIC;
signal DANGLING_U5_r2_11 : STD_LOGIC;
signal DANGLING_U5_r2_10 : STD_LOGIC;
signal DANGLING_U5_r2_9 : STD_LOGIC;
signal DANGLING_U5_r2_8 : STD_LOGIC;
signal DANGLING_U5_r2_7 : STD_LOGIC;
signal DANGLING_U5_r2_6 : STD_LOGIC;
signal DANGLING_U5_r2_5 : STD_LOGIC;
signal DANGLING_U5_r2_4 : STD_LOGIC;
signal DANGLING_U5_r2_3 : STD_LOGIC;
signal DANGLING_U5_r2_2 : STD_LOGIC;
signal DANGLING_U5_r2_1 : STD_LOGIC;
signal DANGLING_U5_r2_0 : STD_LOGIC;
signal DANGLING_U5_r3_126 : STD_LOGIC;
signal DANGLING_U5_r3_125 : STD_LOGIC;
signal DANGLING_U5_r3_124 : STD_LOGIC;
signal DANGLING_U5_r3_123 : STD_LOGIC;
signal DANGLING_U5_r3_122 : STD_LOGIC;
signal DANGLING_U5_r3_121 : STD_LOGIC;
signal DANGLING_U5_r3_120 : STD_LOGIC;
signal DANGLING_U5_r3_119 : STD_LOGIC;
signal DANGLING_U5_r3_118 : STD_LOGIC;
signal DANGLING_U5_r3_117 : STD_LOGIC;
signal DANGLING_U5_r3_116 : STD_LOGIC;
signal DANGLING_U5_r3_115 : STD_LOGIC;
signal DANGLING_U5_r3_114 : STD_LOGIC;
signal DANGLING_U5_r3_113 : STD_LOGIC;
signal DANGLING_U5_r3_112 : STD_LOGIC;
signal DANGLING_U5_r3_111 : STD_LOGIC;
signal DANGLING_U5_r3_110 : STD_LOGIC;
signal DANGLING_U5_r3_109 : STD_LOGIC;
signal DANGLING_U5_r3_108 : STD_LOGIC;
signal DANGLING_U5_r3_107 : STD_LOGIC;
signal DANGLING_U5_r3_106 : STD_LOGIC;
signal DANGLING_U5_r3_105 : STD_LOGIC;
signal DANGLING_U5_r3_104 : STD_LOGIC;
signal DANGLING_U5_r3_103 : STD_LOGIC;
signal DANGLING_U5_r3_102 : STD_LOGIC;
signal DANGLING_U5_r3_101 : STD_LOGIC;
signal DANGLING_U5_r3_100 : STD_LOGIC;
signal DANGLING_U5_r3_99 : STD_LOGIC;
signal DANGLING_U5_r3_98 : STD_LOGIC;
signal DANGLING_U5_r3_97 : STD_LOGIC;
signal DANGLING_U5_r3_96 : STD_LOGIC;
signal DANGLING_U5_r3_95 : STD_LOGIC;
signal DANGLING_U5_r3_94 : STD_LOGIC;
signal DANGLING_U5_r3_93 : STD_LOGIC;
signal DANGLING_U5_r3_92 : STD_LOGIC;
signal DANGLING_U5_r3_91 : STD_LOGIC;
signal DANGLING_U5_r3_90 : STD_LOGIC;
signal DANGLING_U5_r3_89 : STD_LOGIC;
signal DANGLING_U5_r3_88 : STD_LOGIC;
signal DANGLING_U5_r3_87 : STD_LOGIC;
signal DANGLING_U5_r3_86 : STD_LOGIC;
signal DANGLING_U5_r3_85 : STD_LOGIC;
signal DANGLING_U5_r3_84 : STD_LOGIC;
signal DANGLING_U5_r3_83 : STD_LOGIC;
signal DANGLING_U5_r3_82 : STD_LOGIC;
signal DANGLING_U5_r3_81 : STD_LOGIC;
signal DANGLING_U5_r3_80 : STD_LOGIC;
signal DANGLING_U5_r3_79 : STD_LOGIC;
signal DANGLING_U5_r3_78 : STD_LOGIC;
signal DANGLING_U5_r3_77 : STD_LOGIC;
signal DANGLING_U5_r3_76 : STD_LOGIC;
signal DANGLING_U5_r3_75 : STD_LOGIC;
signal DANGLING_U5_r3_74 : STD_LOGIC;
signal DANGLING_U5_r3_73 : STD_LOGIC;
signal DANGLING_U5_r3_72 : STD_LOGIC;
signal DANGLING_U5_r3_71 : STD_LOGIC;
signal DANGLING_U5_r3_70 : STD_LOGIC;
signal DANGLING_U5_r3_69 : STD_LOGIC;
signal DANGLING_U5_r3_68 : STD_LOGIC;
signal DANGLING_U5_r3_67 : STD_LOGIC;
signal DANGLING_U5_r3_66 : STD_LOGIC;
signal DANGLING_U5_r3_65 : STD_LOGIC;
signal DANGLING_U5_r3_64 : STD_LOGIC;
signal DANGLING_U5_r3_63 : STD_LOGIC;
signal DANGLING_U5_r3_62 : STD_LOGIC;
signal DANGLING_U5_r3_61 : STD_LOGIC;
signal DANGLING_U5_r3_60 : STD_LOGIC;
signal DANGLING_U5_r3_59 : STD_LOGIC;
signal DANGLING_U5_r3_58 : STD_LOGIC;
signal DANGLING_U5_r3_57 : STD_LOGIC;
signal DANGLING_U5_r3_56 : STD_LOGIC;
signal DANGLING_U5_r3_55 : STD_LOGIC;
signal DANGLING_U5_r3_54 : STD_LOGIC;
signal DANGLING_U5_r3_53 : STD_LOGIC;
signal DANGLING_U5_r3_52 : STD_LOGIC;
signal DANGLING_U5_r3_51 : STD_LOGIC;
signal DANGLING_U5_r3_50 : STD_LOGIC;
signal DANGLING_U5_r3_49 : STD_LOGIC;
signal DANGLING_U5_r3_48 : STD_LOGIC;
signal DANGLING_U5_r3_47 : STD_LOGIC;
signal DANGLING_U5_r3_46 : STD_LOGIC;
signal DANGLING_U5_r3_45 : STD_LOGIC;
signal DANGLING_U5_r3_44 : STD_LOGIC;
signal DANGLING_U5_r3_43 : STD_LOGIC;
signal DANGLING_U5_r3_42 : STD_LOGIC;
signal DANGLING_U5_r3_41 : STD_LOGIC;
signal DANGLING_U5_r3_40 : STD_LOGIC;
signal DANGLING_U5_r3_39 : STD_LOGIC;
signal DANGLING_U5_r3_38 : STD_LOGIC;
signal DANGLING_U5_r3_37 : STD_LOGIC;
signal DANGLING_U5_r3_36 : STD_LOGIC;
signal DANGLING_U5_r3_35 : STD_LOGIC;
signal DANGLING_U5_r3_34 : STD_LOGIC;
signal DANGLING_U5_r3_33 : STD_LOGIC;
signal DANGLING_U5_r3_32 : STD_LOGIC;
signal DANGLING_U5_r3_31 : STD_LOGIC;
signal DANGLING_U5_r3_30 : STD_LOGIC;
signal DANGLING_U5_r3_29 : STD_LOGIC;
signal DANGLING_U5_r3_28 : STD_LOGIC;
signal DANGLING_U5_r3_27 : STD_LOGIC;
signal DANGLING_U5_r3_26 : STD_LOGIC;
signal DANGLING_U5_r3_25 : STD_LOGIC;
signal DANGLING_U5_r3_24 : STD_LOGIC;
signal DANGLING_U5_r3_23 : STD_LOGIC;
signal DANGLING_U5_r3_22 : STD_LOGIC;
signal DANGLING_U5_r3_21 : STD_LOGIC;
signal DANGLING_U5_r3_20 : STD_LOGIC;
signal DANGLING_U5_r3_19 : STD_LOGIC;
signal DANGLING_U5_r3_18 : STD_LOGIC;
signal DANGLING_U5_r3_17 : STD_LOGIC;
signal DANGLING_U5_r3_16 : STD_LOGIC;
signal DANGLING_U5_r3_15 : STD_LOGIC;
signal DANGLING_U5_r3_14 : STD_LOGIC;
signal DANGLING_U5_r3_13 : STD_LOGIC;
signal DANGLING_U5_r3_12 : STD_LOGIC;
signal DANGLING_U5_r3_11 : STD_LOGIC;
signal DANGLING_U5_r3_10 : STD_LOGIC;
signal DANGLING_U5_r3_9 : STD_LOGIC;
signal DANGLING_U5_r3_8 : STD_LOGIC;
signal DANGLING_U5_r3_7 : STD_LOGIC;
signal DANGLING_U5_r3_6 : STD_LOGIC;
signal DANGLING_U5_r3_5 : STD_LOGIC;
signal DANGLING_U5_r3_4 : STD_LOGIC;
signal DANGLING_U5_r3_3 : STD_LOGIC;
signal DANGLING_U5_r3_2 : STD_LOGIC;
signal DANGLING_U5_r3_1 : STD_LOGIC;
signal DANGLING_U5_r3_0 : STD_LOGIC;
signal DANGLING_U5_ins_out_23 : STD_LOGIC;
signal DANGLING_U5_ins_out_22 : STD_LOGIC;
signal DANGLING_U5_ins_out_21 : STD_LOGIC;
signal DANGLING_U5_ins_out_20 : STD_LOGIC;
signal DANGLING_U5_ins_out_19 : STD_LOGIC;
signal DANGLING_U5_ins_out_18 : STD_LOGIC;
signal DANGLING_U5_ins_out_17 : STD_LOGIC;
signal DANGLING_U5_ins_out_16 : STD_LOGIC;
signal DANGLING_U5_ins_out_15 : STD_LOGIC;
signal DANGLING_U5_ins_out_14 : STD_LOGIC;
signal DANGLING_U5_ins_out_13 : STD_LOGIC;
signal DANGLING_U5_ins_out_12 : STD_LOGIC;
signal DANGLING_U5_ins_out_11 : STD_LOGIC;
signal DANGLING_U5_ins_out_10 : STD_LOGIC;
signal DANGLING_U5_ins_out_9 : STD_LOGIC;
signal DANGLING_U5_ins_out_8 : STD_LOGIC;
signal DANGLING_U5_ins_out_7 : STD_LOGIC;
signal DANGLING_U5_ins_out_6 : STD_LOGIC;
signal DANGLING_U5_ins_out_5 : STD_LOGIC;
signal DANGLING_U5_ins_out_4 : STD_LOGIC;
signal DANGLING_U5_ins_out_3 : STD_LOGIC;
signal DANGLING_U5_ins_out_2 : STD_LOGIC;
signal DANGLING_U5_ins_out_1 : STD_LOGIC;
signal DANGLING_U5_ins_out_0 : STD_LOGIC;

begin

----  Component instantiations  ----

U1 : ins_buffer
  port map(
       ins_out(0) => DANGLING_U1_ins_out_0,
       ins_out(1) => DANGLING_U1_ins_out_1,
       ins_out(2) => DANGLING_U1_ins_out_2,
       ins_out(3) => DANGLING_U1_ins_out_3,
       ins_out(4) => DANGLING_U1_ins_out_4,
       ins_out(5) => DANGLING_U1_ins_out_5,
       ins_out(6) => DANGLING_U1_ins_out_6,
       ins_out(7) => DANGLING_U1_ins_out_7,
       ins_out(8) => DANGLING_U1_ins_out_8,
       ins_out(9) => DANGLING_U1_ins_out_9,
       ins_out(10) => DANGLING_U1_ins_out_10,
       ins_out(11) => DANGLING_U1_ins_out_11,
       ins_out(12) => DANGLING_U1_ins_out_12,
       ins_out(13) => DANGLING_U1_ins_out_13,
       ins_out(14) => DANGLING_U1_ins_out_14,
       ins_out(15) => DANGLING_U1_ins_out_15,
       ins_out(16) => DANGLING_U1_ins_out_16,
       ins_out(17) => DANGLING_U1_ins_out_17,
       ins_out(18) => DANGLING_U1_ins_out_18,
       ins_out(19) => DANGLING_U1_ins_out_19,
       ins_out(20) => DANGLING_U1_ins_out_20,
       ins_out(21) => DANGLING_U1_ins_out_21,
       ins_out(22) => DANGLING_U1_ins_out_22,
       ins_out(23) => DANGLING_U1_ins_out_23,
       ins_out(24) => NET114,
       clk => clk,
       instructions => instruction
  );

U2 : alu
  port map(
       alu_out(0) => DANGLING_U2_alu_out_0,
       alu_out(1) => DANGLING_U2_alu_out_1,
       alu_out(2) => DANGLING_U2_alu_out_2,
       alu_out(3) => DANGLING_U2_alu_out_3,
       alu_out(4) => DANGLING_U2_alu_out_4,
       alu_out(5) => DANGLING_U2_alu_out_5,
       alu_out(6) => DANGLING_U2_alu_out_6,
       alu_out(7) => DANGLING_U2_alu_out_7,
       alu_out(8) => DANGLING_U2_alu_out_8,
       alu_out(9) => DANGLING_U2_alu_out_9,
       alu_out(10) => DANGLING_U2_alu_out_10,
       alu_out(11) => DANGLING_U2_alu_out_11,
       alu_out(12) => DANGLING_U2_alu_out_12,
       alu_out(13) => DANGLING_U2_alu_out_13,
       alu_out(14) => DANGLING_U2_alu_out_14,
       alu_out(15) => DANGLING_U2_alu_out_15,
       alu_out(16) => DANGLING_U2_alu_out_16,
       alu_out(17) => DANGLING_U2_alu_out_17,
       alu_out(18) => DANGLING_U2_alu_out_18,
       alu_out(19) => DANGLING_U2_alu_out_19,
       alu_out(20) => DANGLING_U2_alu_out_20,
       alu_out(21) => DANGLING_U2_alu_out_21,
       alu_out(22) => DANGLING_U2_alu_out_22,
       alu_out(23) => DANGLING_U2_alu_out_23,
       alu_out(24) => DANGLING_U2_alu_out_24,
       alu_out(25) => DANGLING_U2_alu_out_25,
       alu_out(26) => DANGLING_U2_alu_out_26,
       alu_out(27) => DANGLING_U2_alu_out_27,
       alu_out(28) => DANGLING_U2_alu_out_28,
       alu_out(29) => DANGLING_U2_alu_out_29,
       alu_out(30) => DANGLING_U2_alu_out_30,
       alu_out(31) => DANGLING_U2_alu_out_31,
       alu_out(32) => DANGLING_U2_alu_out_32,
       alu_out(33) => DANGLING_U2_alu_out_33,
       alu_out(34) => DANGLING_U2_alu_out_34,
       alu_out(35) => DANGLING_U2_alu_out_35,
       alu_out(36) => DANGLING_U2_alu_out_36,
       alu_out(37) => DANGLING_U2_alu_out_37,
       alu_out(38) => DANGLING_U2_alu_out_38,
       alu_out(39) => DANGLING_U2_alu_out_39,
       alu_out(40) => DANGLING_U2_alu_out_40,
       alu_out(41) => DANGLING_U2_alu_out_41,
       alu_out(42) => DANGLING_U2_alu_out_42,
       alu_out(43) => DANGLING_U2_alu_out_43,
       alu_out(44) => DANGLING_U2_alu_out_44,
       alu_out(45) => DANGLING_U2_alu_out_45,
       alu_out(46) => DANGLING_U2_alu_out_46,
       alu_out(47) => DANGLING_U2_alu_out_47,
       alu_out(48) => DANGLING_U2_alu_out_48,
       alu_out(49) => DANGLING_U2_alu_out_49,
       alu_out(50) => DANGLING_U2_alu_out_50,
       alu_out(51) => DANGLING_U2_alu_out_51,
       alu_out(52) => DANGLING_U2_alu_out_52,
       alu_out(53) => DANGLING_U2_alu_out_53,
       alu_out(54) => DANGLING_U2_alu_out_54,
       alu_out(55) => DANGLING_U2_alu_out_55,
       alu_out(56) => DANGLING_U2_alu_out_56,
       alu_out(57) => DANGLING_U2_alu_out_57,
       alu_out(58) => DANGLING_U2_alu_out_58,
       alu_out(59) => DANGLING_U2_alu_out_59,
       alu_out(60) => DANGLING_U2_alu_out_60,
       alu_out(61) => DANGLING_U2_alu_out_61,
       alu_out(62) => DANGLING_U2_alu_out_62,
       alu_out(63) => DANGLING_U2_alu_out_63,
       alu_out(64) => DANGLING_U2_alu_out_64,
       alu_out(65) => DANGLING_U2_alu_out_65,
       alu_out(66) => DANGLING_U2_alu_out_66,
       alu_out(67) => DANGLING_U2_alu_out_67,
       alu_out(68) => DANGLING_U2_alu_out_68,
       alu_out(69) => DANGLING_U2_alu_out_69,
       alu_out(70) => DANGLING_U2_alu_out_70,
       alu_out(71) => DANGLING_U2_alu_out_71,
       alu_out(72) => DANGLING_U2_alu_out_72,
       alu_out(73) => DANGLING_U2_alu_out_73,
       alu_out(74) => DANGLING_U2_alu_out_74,
       alu_out(75) => DANGLING_U2_alu_out_75,
       alu_out(76) => DANGLING_U2_alu_out_76,
       alu_out(77) => DANGLING_U2_alu_out_77,
       alu_out(78) => DANGLING_U2_alu_out_78,
       alu_out(79) => DANGLING_U2_alu_out_79,
       alu_out(80) => DANGLING_U2_alu_out_80,
       alu_out(81) => DANGLING_U2_alu_out_81,
       alu_out(82) => DANGLING_U2_alu_out_82,
       alu_out(83) => DANGLING_U2_alu_out_83,
       alu_out(84) => DANGLING_U2_alu_out_84,
       alu_out(85) => DANGLING_U2_alu_out_85,
       alu_out(86) => DANGLING_U2_alu_out_86,
       alu_out(87) => DANGLING_U2_alu_out_87,
       alu_out(88) => DANGLING_U2_alu_out_88,
       alu_out(89) => DANGLING_U2_alu_out_89,
       alu_out(90) => DANGLING_U2_alu_out_90,
       alu_out(91) => DANGLING_U2_alu_out_91,
       alu_out(92) => DANGLING_U2_alu_out_92,
       alu_out(93) => DANGLING_U2_alu_out_93,
       alu_out(94) => DANGLING_U2_alu_out_94,
       alu_out(95) => DANGLING_U2_alu_out_95,
       alu_out(96) => DANGLING_U2_alu_out_96,
       alu_out(97) => DANGLING_U2_alu_out_97,
       alu_out(98) => DANGLING_U2_alu_out_98,
       alu_out(99) => DANGLING_U2_alu_out_99,
       alu_out(100) => DANGLING_U2_alu_out_100,
       alu_out(101) => DANGLING_U2_alu_out_101,
       alu_out(102) => DANGLING_U2_alu_out_102,
       alu_out(103) => DANGLING_U2_alu_out_103,
       alu_out(104) => DANGLING_U2_alu_out_104,
       alu_out(105) => DANGLING_U2_alu_out_105,
       alu_out(106) => DANGLING_U2_alu_out_106,
       alu_out(107) => DANGLING_U2_alu_out_107,
       alu_out(108) => DANGLING_U2_alu_out_108,
       alu_out(109) => DANGLING_U2_alu_out_109,
       alu_out(110) => DANGLING_U2_alu_out_110,
       alu_out(111) => DANGLING_U2_alu_out_111,
       alu_out(112) => DANGLING_U2_alu_out_112,
       alu_out(113) => DANGLING_U2_alu_out_113,
       alu_out(114) => DANGLING_U2_alu_out_114,
       alu_out(115) => DANGLING_U2_alu_out_115,
       alu_out(116) => DANGLING_U2_alu_out_116,
       alu_out(117) => DANGLING_U2_alu_out_117,
       alu_out(118) => DANGLING_U2_alu_out_118,
       alu_out(119) => DANGLING_U2_alu_out_119,
       alu_out(120) => DANGLING_U2_alu_out_120,
       alu_out(121) => DANGLING_U2_alu_out_121,
       alu_out(122) => DANGLING_U2_alu_out_122,
       alu_out(123) => DANGLING_U2_alu_out_123,
       alu_out(124) => DANGLING_U2_alu_out_124,
       alu_out(125) => DANGLING_U2_alu_out_125,
       alu_out(126) => DANGLING_U2_alu_out_126,
       alu_out(127) => NET210,
       ins(0) => Dangling_Input_Signal,
       ins(1) => Dangling_Input_Signal,
       ins(2) => Dangling_Input_Signal,
       ins(3) => Dangling_Input_Signal,
       ins(4) => Dangling_Input_Signal,
       ins(5) => Dangling_Input_Signal,
       ins(6) => Dangling_Input_Signal,
       ins(7) => Dangling_Input_Signal,
       ins(8) => Dangling_Input_Signal,
       ins(9) => Dangling_Input_Signal,
       ins(10) => Dangling_Input_Signal,
       ins(11) => Dangling_Input_Signal,
       ins(12) => Dangling_Input_Signal,
       ins(13) => Dangling_Input_Signal,
       ins(14) => Dangling_Input_Signal,
       ins(15) => Dangling_Input_Signal,
       ins(16) => Dangling_Input_Signal,
       ins(17) => Dangling_Input_Signal,
       ins(18) => Dangling_Input_Signal,
       ins(19) => Dangling_Input_Signal,
       ins(20) => Dangling_Input_Signal,
       ins(21) => Dangling_Input_Signal,
       ins(22) => Dangling_Input_Signal,
       ins(23) => Dangling_Input_Signal,
       ins(24) => Dangling_Input_Signal,
       ins_out(0) => DANGLING_U2_ins_out_0,
       ins_out(1) => DANGLING_U2_ins_out_1,
       ins_out(2) => DANGLING_U2_ins_out_2,
       ins_out(3) => DANGLING_U2_ins_out_3,
       ins_out(4) => DANGLING_U2_ins_out_4,
       ins_out(5) => DANGLING_U2_ins_out_5,
       ins_out(6) => DANGLING_U2_ins_out_6,
       ins_out(7) => DANGLING_U2_ins_out_7,
       ins_out(8) => DANGLING_U2_ins_out_8,
       ins_out(9) => DANGLING_U2_ins_out_9,
       ins_out(10) => DANGLING_U2_ins_out_10,
       ins_out(11) => DANGLING_U2_ins_out_11,
       ins_out(12) => DANGLING_U2_ins_out_12,
       ins_out(13) => DANGLING_U2_ins_out_13,
       ins_out(14) => DANGLING_U2_ins_out_14,
       ins_out(15) => DANGLING_U2_ins_out_15,
       ins_out(16) => DANGLING_U2_ins_out_16,
       ins_out(17) => DANGLING_U2_ins_out_17,
       ins_out(18) => DANGLING_U2_ins_out_18,
       ins_out(19) => DANGLING_U2_ins_out_19,
       ins_out(20) => DANGLING_U2_ins_out_20,
       ins_out(21) => DANGLING_U2_ins_out_21,
       ins_out(22) => DANGLING_U2_ins_out_22,
       ins_out(23) => DANGLING_U2_ins_out_23,
       ins_out(24) => NET246,
       r1(0) => Dangling_Input_Signal,
       r1(1) => Dangling_Input_Signal,
       r1(2) => Dangling_Input_Signal,
       r1(3) => Dangling_Input_Signal,
       r1(4) => Dangling_Input_Signal,
       r1(5) => Dangling_Input_Signal,
       r1(6) => Dangling_Input_Signal,
       r1(7) => Dangling_Input_Signal,
       r1(8) => Dangling_Input_Signal,
       r1(9) => Dangling_Input_Signal,
       r1(10) => Dangling_Input_Signal,
       r1(11) => Dangling_Input_Signal,
       r1(12) => Dangling_Input_Signal,
       r1(13) => Dangling_Input_Signal,
       r1(14) => Dangling_Input_Signal,
       r1(15) => Dangling_Input_Signal,
       r1(16) => Dangling_Input_Signal,
       r1(17) => Dangling_Input_Signal,
       r1(18) => Dangling_Input_Signal,
       r1(19) => Dangling_Input_Signal,
       r1(20) => Dangling_Input_Signal,
       r1(21) => Dangling_Input_Signal,
       r1(22) => Dangling_Input_Signal,
       r1(23) => Dangling_Input_Signal,
       r1(24) => Dangling_Input_Signal,
       r1(25) => Dangling_Input_Signal,
       r1(26) => Dangling_Input_Signal,
       r1(27) => Dangling_Input_Signal,
       r1(28) => Dangling_Input_Signal,
       r1(29) => Dangling_Input_Signal,
       r1(30) => Dangling_Input_Signal,
       r1(31) => Dangling_Input_Signal,
       r1(32) => Dangling_Input_Signal,
       r1(33) => Dangling_Input_Signal,
       r1(34) => Dangling_Input_Signal,
       r1(35) => Dangling_Input_Signal,
       r1(36) => Dangling_Input_Signal,
       r1(37) => Dangling_Input_Signal,
       r1(38) => Dangling_Input_Signal,
       r1(39) => Dangling_Input_Signal,
       r1(40) => Dangling_Input_Signal,
       r1(41) => Dangling_Input_Signal,
       r1(42) => Dangling_Input_Signal,
       r1(43) => Dangling_Input_Signal,
       r1(44) => Dangling_Input_Signal,
       r1(45) => Dangling_Input_Signal,
       r1(46) => Dangling_Input_Signal,
       r1(47) => Dangling_Input_Signal,
       r1(48) => Dangling_Input_Signal,
       r1(49) => Dangling_Input_Signal,
       r1(50) => Dangling_Input_Signal,
       r1(51) => Dangling_Input_Signal,
       r1(52) => Dangling_Input_Signal,
       r1(53) => Dangling_Input_Signal,
       r1(54) => Dangling_Input_Signal,
       r1(55) => Dangling_Input_Signal,
       r1(56) => Dangling_Input_Signal,
       r1(57) => Dangling_Input_Signal,
       r1(58) => Dangling_Input_Signal,
       r1(59) => Dangling_Input_Signal,
       r1(60) => Dangling_Input_Signal,
       r1(61) => Dangling_Input_Signal,
       r1(62) => Dangling_Input_Signal,
       r1(63) => Dangling_Input_Signal,
       r1(64) => Dangling_Input_Signal,
       r1(65) => Dangling_Input_Signal,
       r1(66) => Dangling_Input_Signal,
       r1(67) => Dangling_Input_Signal,
       r1(68) => Dangling_Input_Signal,
       r1(69) => Dangling_Input_Signal,
       r1(70) => Dangling_Input_Signal,
       r1(71) => Dangling_Input_Signal,
       r1(72) => Dangling_Input_Signal,
       r1(73) => Dangling_Input_Signal,
       r1(74) => Dangling_Input_Signal,
       r1(75) => Dangling_Input_Signal,
       r1(76) => Dangling_Input_Signal,
       r1(77) => Dangling_Input_Signal,
       r1(78) => Dangling_Input_Signal,
       r1(79) => Dangling_Input_Signal,
       r1(80) => Dangling_Input_Signal,
       r1(81) => Dangling_Input_Signal,
       r1(82) => Dangling_Input_Signal,
       r1(83) => Dangling_Input_Signal,
       r1(84) => Dangling_Input_Signal,
       r1(85) => Dangling_Input_Signal,
       r1(86) => Dangling_Input_Signal,
       r1(87) => Dangling_Input_Signal,
       r1(88) => Dangling_Input_Signal,
       r1(89) => Dangling_Input_Signal,
       r1(90) => Dangling_Input_Signal,
       r1(91) => Dangling_Input_Signal,
       r1(92) => Dangling_Input_Signal,
       r1(93) => Dangling_Input_Signal,
       r1(94) => Dangling_Input_Signal,
       r1(95) => Dangling_Input_Signal,
       r1(96) => Dangling_Input_Signal,
       r1(97) => Dangling_Input_Signal,
       r1(98) => Dangling_Input_Signal,
       r1(99) => Dangling_Input_Signal,
       r1(100) => Dangling_Input_Signal,
       r1(101) => Dangling_Input_Signal,
       r1(102) => Dangling_Input_Signal,
       r1(103) => Dangling_Input_Signal,
       r1(104) => Dangling_Input_Signal,
       r1(105) => Dangling_Input_Signal,
       r1(106) => Dangling_Input_Signal,
       r1(107) => Dangling_Input_Signal,
       r1(108) => Dangling_Input_Signal,
       r1(109) => Dangling_Input_Signal,
       r1(110) => Dangling_Input_Signal,
       r1(111) => Dangling_Input_Signal,
       r1(112) => Dangling_Input_Signal,
       r1(113) => Dangling_Input_Signal,
       r1(114) => Dangling_Input_Signal,
       r1(115) => Dangling_Input_Signal,
       r1(116) => Dangling_Input_Signal,
       r1(117) => Dangling_Input_Signal,
       r1(118) => Dangling_Input_Signal,
       r1(119) => Dangling_Input_Signal,
       r1(120) => Dangling_Input_Signal,
       r1(121) => Dangling_Input_Signal,
       r1(122) => Dangling_Input_Signal,
       r1(123) => Dangling_Input_Signal,
       r1(124) => Dangling_Input_Signal,
       r1(125) => Dangling_Input_Signal,
       r1(126) => Dangling_Input_Signal,
       r1(127) => NET238,
       r2(0) => Dangling_Input_Signal,
       r2(1) => Dangling_Input_Signal,
       r2(2) => Dangling_Input_Signal,
       r2(3) => Dangling_Input_Signal,
       r2(4) => Dangling_Input_Signal,
       r2(5) => Dangling_Input_Signal,
       r2(6) => Dangling_Input_Signal,
       r2(7) => Dangling_Input_Signal,
       r2(8) => Dangling_Input_Signal,
       r2(9) => Dangling_Input_Signal,
       r2(10) => Dangling_Input_Signal,
       r2(11) => Dangling_Input_Signal,
       r2(12) => Dangling_Input_Signal,
       r2(13) => Dangling_Input_Signal,
       r2(14) => Dangling_Input_Signal,
       r2(15) => Dangling_Input_Signal,
       r2(16) => Dangling_Input_Signal,
       r2(17) => Dangling_Input_Signal,
       r2(18) => Dangling_Input_Signal,
       r2(19) => Dangling_Input_Signal,
       r2(20) => Dangling_Input_Signal,
       r2(21) => Dangling_Input_Signal,
       r2(22) => Dangling_Input_Signal,
       r2(23) => Dangling_Input_Signal,
       r2(24) => Dangling_Input_Signal,
       r2(25) => Dangling_Input_Signal,
       r2(26) => Dangling_Input_Signal,
       r2(27) => Dangling_Input_Signal,
       r2(28) => Dangling_Input_Signal,
       r2(29) => Dangling_Input_Signal,
       r2(30) => Dangling_Input_Signal,
       r2(31) => Dangling_Input_Signal,
       r2(32) => Dangling_Input_Signal,
       r2(33) => Dangling_Input_Signal,
       r2(34) => Dangling_Input_Signal,
       r2(35) => Dangling_Input_Signal,
       r2(36) => Dangling_Input_Signal,
       r2(37) => Dangling_Input_Signal,
       r2(38) => Dangling_Input_Signal,
       r2(39) => Dangling_Input_Signal,
       r2(40) => Dangling_Input_Signal,
       r2(41) => Dangling_Input_Signal,
       r2(42) => Dangling_Input_Signal,
       r2(43) => Dangling_Input_Signal,
       r2(44) => Dangling_Input_Signal,
       r2(45) => Dangling_Input_Signal,
       r2(46) => Dangling_Input_Signal,
       r2(47) => Dangling_Input_Signal,
       r2(48) => Dangling_Input_Signal,
       r2(49) => Dangling_Input_Signal,
       r2(50) => Dangling_Input_Signal,
       r2(51) => Dangling_Input_Signal,
       r2(52) => Dangling_Input_Signal,
       r2(53) => Dangling_Input_Signal,
       r2(54) => Dangling_Input_Signal,
       r2(55) => Dangling_Input_Signal,
       r2(56) => Dangling_Input_Signal,
       r2(57) => Dangling_Input_Signal,
       r2(58) => Dangling_Input_Signal,
       r2(59) => Dangling_Input_Signal,
       r2(60) => Dangling_Input_Signal,
       r2(61) => Dangling_Input_Signal,
       r2(62) => Dangling_Input_Signal,
       r2(63) => Dangling_Input_Signal,
       r2(64) => Dangling_Input_Signal,
       r2(65) => Dangling_Input_Signal,
       r2(66) => Dangling_Input_Signal,
       r2(67) => Dangling_Input_Signal,
       r2(68) => Dangling_Input_Signal,
       r2(69) => Dangling_Input_Signal,
       r2(70) => Dangling_Input_Signal,
       r2(71) => Dangling_Input_Signal,
       r2(72) => Dangling_Input_Signal,
       r2(73) => Dangling_Input_Signal,
       r2(74) => Dangling_Input_Signal,
       r2(75) => Dangling_Input_Signal,
       r2(76) => Dangling_Input_Signal,
       r2(77) => Dangling_Input_Signal,
       r2(78) => Dangling_Input_Signal,
       r2(79) => Dangling_Input_Signal,
       r2(80) => Dangling_Input_Signal,
       r2(81) => Dangling_Input_Signal,
       r2(82) => Dangling_Input_Signal,
       r2(83) => Dangling_Input_Signal,
       r2(84) => Dangling_Input_Signal,
       r2(85) => Dangling_Input_Signal,
       r2(86) => Dangling_Input_Signal,
       r2(87) => Dangling_Input_Signal,
       r2(88) => Dangling_Input_Signal,
       r2(89) => Dangling_Input_Signal,
       r2(90) => Dangling_Input_Signal,
       r2(91) => Dangling_Input_Signal,
       r2(92) => Dangling_Input_Signal,
       r2(93) => Dangling_Input_Signal,
       r2(94) => Dangling_Input_Signal,
       r2(95) => Dangling_Input_Signal,
       r2(96) => Dangling_Input_Signal,
       r2(97) => Dangling_Input_Signal,
       r2(98) => Dangling_Input_Signal,
       r2(99) => Dangling_Input_Signal,
       r2(100) => Dangling_Input_Signal,
       r2(101) => Dangling_Input_Signal,
       r2(102) => Dangling_Input_Signal,
       r2(103) => Dangling_Input_Signal,
       r2(104) => Dangling_Input_Signal,
       r2(105) => Dangling_Input_Signal,
       r2(106) => Dangling_Input_Signal,
       r2(107) => Dangling_Input_Signal,
       r2(108) => Dangling_Input_Signal,
       r2(109) => Dangling_Input_Signal,
       r2(110) => Dangling_Input_Signal,
       r2(111) => Dangling_Input_Signal,
       r2(112) => Dangling_Input_Signal,
       r2(113) => Dangling_Input_Signal,
       r2(114) => Dangling_Input_Signal,
       r2(115) => Dangling_Input_Signal,
       r2(116) => Dangling_Input_Signal,
       r2(117) => Dangling_Input_Signal,
       r2(118) => Dangling_Input_Signal,
       r2(119) => Dangling_Input_Signal,
       r2(120) => Dangling_Input_Signal,
       r2(121) => Dangling_Input_Signal,
       r2(122) => Dangling_Input_Signal,
       r2(123) => Dangling_Input_Signal,
       r2(124) => Dangling_Input_Signal,
       r2(125) => Dangling_Input_Signal,
       r2(126) => Dangling_Input_Signal,
       r2(127) => NET230,
       r3(0) => Dangling_Input_Signal,
       r3(1) => Dangling_Input_Signal,
       r3(2) => Dangling_Input_Signal,
       r3(3) => Dangling_Input_Signal,
       r3(4) => Dangling_Input_Signal,
       r3(5) => Dangling_Input_Signal,
       r3(6) => Dangling_Input_Signal,
       r3(7) => Dangling_Input_Signal,
       r3(8) => Dangling_Input_Signal,
       r3(9) => Dangling_Input_Signal,
       r3(10) => Dangling_Input_Signal,
       r3(11) => Dangling_Input_Signal,
       r3(12) => Dangling_Input_Signal,
       r3(13) => Dangling_Input_Signal,
       r3(14) => Dangling_Input_Signal,
       r3(15) => Dangling_Input_Signal,
       r3(16) => Dangling_Input_Signal,
       r3(17) => Dangling_Input_Signal,
       r3(18) => Dangling_Input_Signal,
       r3(19) => Dangling_Input_Signal,
       r3(20) => Dangling_Input_Signal,
       r3(21) => Dangling_Input_Signal,
       r3(22) => Dangling_Input_Signal,
       r3(23) => Dangling_Input_Signal,
       r3(24) => Dangling_Input_Signal,
       r3(25) => Dangling_Input_Signal,
       r3(26) => Dangling_Input_Signal,
       r3(27) => Dangling_Input_Signal,
       r3(28) => Dangling_Input_Signal,
       r3(29) => Dangling_Input_Signal,
       r3(30) => Dangling_Input_Signal,
       r3(31) => Dangling_Input_Signal,
       r3(32) => Dangling_Input_Signal,
       r3(33) => Dangling_Input_Signal,
       r3(34) => Dangling_Input_Signal,
       r3(35) => Dangling_Input_Signal,
       r3(36) => Dangling_Input_Signal,
       r3(37) => Dangling_Input_Signal,
       r3(38) => Dangling_Input_Signal,
       r3(39) => Dangling_Input_Signal,
       r3(40) => Dangling_Input_Signal,
       r3(41) => Dangling_Input_Signal,
       r3(42) => Dangling_Input_Signal,
       r3(43) => Dangling_Input_Signal,
       r3(44) => Dangling_Input_Signal,
       r3(45) => Dangling_Input_Signal,
       r3(46) => Dangling_Input_Signal,
       r3(47) => Dangling_Input_Signal,
       r3(48) => Dangling_Input_Signal,
       r3(49) => Dangling_Input_Signal,
       r3(50) => Dangling_Input_Signal,
       r3(51) => Dangling_Input_Signal,
       r3(52) => Dangling_Input_Signal,
       r3(53) => Dangling_Input_Signal,
       r3(54) => Dangling_Input_Signal,
       r3(55) => Dangling_Input_Signal,
       r3(56) => Dangling_Input_Signal,
       r3(57) => Dangling_Input_Signal,
       r3(58) => Dangling_Input_Signal,
       r3(59) => Dangling_Input_Signal,
       r3(60) => Dangling_Input_Signal,
       r3(61) => Dangling_Input_Signal,
       r3(62) => Dangling_Input_Signal,
       r3(63) => Dangling_Input_Signal,
       r3(64) => Dangling_Input_Signal,
       r3(65) => Dangling_Input_Signal,
       r3(66) => Dangling_Input_Signal,
       r3(67) => Dangling_Input_Signal,
       r3(68) => Dangling_Input_Signal,
       r3(69) => Dangling_Input_Signal,
       r3(70) => Dangling_Input_Signal,
       r3(71) => Dangling_Input_Signal,
       r3(72) => Dangling_Input_Signal,
       r3(73) => Dangling_Input_Signal,
       r3(74) => Dangling_Input_Signal,
       r3(75) => Dangling_Input_Signal,
       r3(76) => Dangling_Input_Signal,
       r3(77) => Dangling_Input_Signal,
       r3(78) => Dangling_Input_Signal,
       r3(79) => Dangling_Input_Signal,
       r3(80) => Dangling_Input_Signal,
       r3(81) => Dangling_Input_Signal,
       r3(82) => Dangling_Input_Signal,
       r3(83) => Dangling_Input_Signal,
       r3(84) => Dangling_Input_Signal,
       r3(85) => Dangling_Input_Signal,
       r3(86) => Dangling_Input_Signal,
       r3(87) => Dangling_Input_Signal,
       r3(88) => Dangling_Input_Signal,
       r3(89) => Dangling_Input_Signal,
       r3(90) => Dangling_Input_Signal,
       r3(91) => Dangling_Input_Signal,
       r3(92) => Dangling_Input_Signal,
       r3(93) => Dangling_Input_Signal,
       r3(94) => Dangling_Input_Signal,
       r3(95) => Dangling_Input_Signal,
       r3(96) => Dangling_Input_Signal,
       r3(97) => Dangling_Input_Signal,
       r3(98) => Dangling_Input_Signal,
       r3(99) => Dangling_Input_Signal,
       r3(100) => Dangling_Input_Signal,
       r3(101) => Dangling_Input_Signal,
       r3(102) => Dangling_Input_Signal,
       r3(103) => Dangling_Input_Signal,
       r3(104) => Dangling_Input_Signal,
       r3(105) => Dangling_Input_Signal,
       r3(106) => Dangling_Input_Signal,
       r3(107) => Dangling_Input_Signal,
       r3(108) => Dangling_Input_Signal,
       r3(109) => Dangling_Input_Signal,
       r3(110) => Dangling_Input_Signal,
       r3(111) => Dangling_Input_Signal,
       r3(112) => Dangling_Input_Signal,
       r3(113) => Dangling_Input_Signal,
       r3(114) => Dangling_Input_Signal,
       r3(115) => Dangling_Input_Signal,
       r3(116) => Dangling_Input_Signal,
       r3(117) => Dangling_Input_Signal,
       r3(118) => Dangling_Input_Signal,
       r3(119) => Dangling_Input_Signal,
       r3(120) => Dangling_Input_Signal,
       r3(121) => Dangling_Input_Signal,
       r3(122) => Dangling_Input_Signal,
       r3(123) => Dangling_Input_Signal,
       r3(124) => Dangling_Input_Signal,
       r3(125) => Dangling_Input_Signal,
       r3(126) => Dangling_Input_Signal,
       r3(127) => NET222,
       clk => clk
  );

U3 : forwarding_unit
  port map(
       ALU_out(0) => Dangling_Input_Signal,
       ALU_out(1) => Dangling_Input_Signal,
       ALU_out(2) => Dangling_Input_Signal,
       ALU_out(3) => Dangling_Input_Signal,
       ALU_out(4) => Dangling_Input_Signal,
       ALU_out(5) => Dangling_Input_Signal,
       ALU_out(6) => Dangling_Input_Signal,
       ALU_out(7) => Dangling_Input_Signal,
       ALU_out(8) => Dangling_Input_Signal,
       ALU_out(9) => Dangling_Input_Signal,
       ALU_out(10) => Dangling_Input_Signal,
       ALU_out(11) => Dangling_Input_Signal,
       ALU_out(12) => Dangling_Input_Signal,
       ALU_out(13) => Dangling_Input_Signal,
       ALU_out(14) => Dangling_Input_Signal,
       ALU_out(15) => Dangling_Input_Signal,
       ALU_out(16) => Dangling_Input_Signal,
       ALU_out(17) => Dangling_Input_Signal,
       ALU_out(18) => Dangling_Input_Signal,
       ALU_out(19) => Dangling_Input_Signal,
       ALU_out(20) => Dangling_Input_Signal,
       ALU_out(21) => Dangling_Input_Signal,
       ALU_out(22) => Dangling_Input_Signal,
       ALU_out(23) => Dangling_Input_Signal,
       ALU_out(24) => Dangling_Input_Signal,
       ALU_out(25) => Dangling_Input_Signal,
       ALU_out(26) => Dangling_Input_Signal,
       ALU_out(27) => Dangling_Input_Signal,
       ALU_out(28) => Dangling_Input_Signal,
       ALU_out(29) => Dangling_Input_Signal,
       ALU_out(30) => Dangling_Input_Signal,
       ALU_out(31) => Dangling_Input_Signal,
       ALU_out(32) => Dangling_Input_Signal,
       ALU_out(33) => Dangling_Input_Signal,
       ALU_out(34) => Dangling_Input_Signal,
       ALU_out(35) => Dangling_Input_Signal,
       ALU_out(36) => Dangling_Input_Signal,
       ALU_out(37) => Dangling_Input_Signal,
       ALU_out(38) => Dangling_Input_Signal,
       ALU_out(39) => Dangling_Input_Signal,
       ALU_out(40) => Dangling_Input_Signal,
       ALU_out(41) => Dangling_Input_Signal,
       ALU_out(42) => Dangling_Input_Signal,
       ALU_out(43) => Dangling_Input_Signal,
       ALU_out(44) => Dangling_Input_Signal,
       ALU_out(45) => Dangling_Input_Signal,
       ALU_out(46) => Dangling_Input_Signal,
       ALU_out(47) => Dangling_Input_Signal,
       ALU_out(48) => Dangling_Input_Signal,
       ALU_out(49) => Dangling_Input_Signal,
       ALU_out(50) => Dangling_Input_Signal,
       ALU_out(51) => Dangling_Input_Signal,
       ALU_out(52) => Dangling_Input_Signal,
       ALU_out(53) => Dangling_Input_Signal,
       ALU_out(54) => Dangling_Input_Signal,
       ALU_out(55) => Dangling_Input_Signal,
       ALU_out(56) => Dangling_Input_Signal,
       ALU_out(57) => Dangling_Input_Signal,
       ALU_out(58) => Dangling_Input_Signal,
       ALU_out(59) => Dangling_Input_Signal,
       ALU_out(60) => Dangling_Input_Signal,
       ALU_out(61) => Dangling_Input_Signal,
       ALU_out(62) => Dangling_Input_Signal,
       ALU_out(63) => Dangling_Input_Signal,
       ALU_out(64) => Dangling_Input_Signal,
       ALU_out(65) => Dangling_Input_Signal,
       ALU_out(66) => Dangling_Input_Signal,
       ALU_out(67) => Dangling_Input_Signal,
       ALU_out(68) => Dangling_Input_Signal,
       ALU_out(69) => Dangling_Input_Signal,
       ALU_out(70) => Dangling_Input_Signal,
       ALU_out(71) => Dangling_Input_Signal,
       ALU_out(72) => Dangling_Input_Signal,
       ALU_out(73) => Dangling_Input_Signal,
       ALU_out(74) => Dangling_Input_Signal,
       ALU_out(75) => Dangling_Input_Signal,
       ALU_out(76) => Dangling_Input_Signal,
       ALU_out(77) => Dangling_Input_Signal,
       ALU_out(78) => Dangling_Input_Signal,
       ALU_out(79) => Dangling_Input_Signal,
       ALU_out(80) => Dangling_Input_Signal,
       ALU_out(81) => Dangling_Input_Signal,
       ALU_out(82) => Dangling_Input_Signal,
       ALU_out(83) => Dangling_Input_Signal,
       ALU_out(84) => Dangling_Input_Signal,
       ALU_out(85) => Dangling_Input_Signal,
       ALU_out(86) => Dangling_Input_Signal,
       ALU_out(87) => Dangling_Input_Signal,
       ALU_out(88) => Dangling_Input_Signal,
       ALU_out(89) => Dangling_Input_Signal,
       ALU_out(90) => Dangling_Input_Signal,
       ALU_out(91) => Dangling_Input_Signal,
       ALU_out(92) => Dangling_Input_Signal,
       ALU_out(93) => Dangling_Input_Signal,
       ALU_out(94) => Dangling_Input_Signal,
       ALU_out(95) => Dangling_Input_Signal,
       ALU_out(96) => Dangling_Input_Signal,
       ALU_out(97) => Dangling_Input_Signal,
       ALU_out(98) => Dangling_Input_Signal,
       ALU_out(99) => Dangling_Input_Signal,
       ALU_out(100) => Dangling_Input_Signal,
       ALU_out(101) => Dangling_Input_Signal,
       ALU_out(102) => Dangling_Input_Signal,
       ALU_out(103) => Dangling_Input_Signal,
       ALU_out(104) => Dangling_Input_Signal,
       ALU_out(105) => Dangling_Input_Signal,
       ALU_out(106) => Dangling_Input_Signal,
       ALU_out(107) => Dangling_Input_Signal,
       ALU_out(108) => Dangling_Input_Signal,
       ALU_out(109) => Dangling_Input_Signal,
       ALU_out(110) => Dangling_Input_Signal,
       ALU_out(111) => Dangling_Input_Signal,
       ALU_out(112) => Dangling_Input_Signal,
       ALU_out(113) => Dangling_Input_Signal,
       ALU_out(114) => Dangling_Input_Signal,
       ALU_out(115) => Dangling_Input_Signal,
       ALU_out(116) => Dangling_Input_Signal,
       ALU_out(117) => Dangling_Input_Signal,
       ALU_out(118) => Dangling_Input_Signal,
       ALU_out(119) => Dangling_Input_Signal,
       ALU_out(120) => Dangling_Input_Signal,
       ALU_out(121) => Dangling_Input_Signal,
       ALU_out(122) => Dangling_Input_Signal,
       ALU_out(123) => Dangling_Input_Signal,
       ALU_out(124) => Dangling_Input_Signal,
       ALU_out(125) => Dangling_Input_Signal,
       ALU_out(126) => Dangling_Input_Signal,
       ALU_out(127) => NET210,
       ins(0) => Dangling_Input_Signal,
       ins(1) => Dangling_Input_Signal,
       ins(2) => Dangling_Input_Signal,
       ins(3) => Dangling_Input_Signal,
       ins(4) => Dangling_Input_Signal,
       ins(5) => Dangling_Input_Signal,
       ins(6) => Dangling_Input_Signal,
       ins(7) => Dangling_Input_Signal,
       ins(8) => Dangling_Input_Signal,
       ins(9) => Dangling_Input_Signal,
       ins(10) => Dangling_Input_Signal,
       ins(11) => Dangling_Input_Signal,
       ins(12) => Dangling_Input_Signal,
       ins(13) => Dangling_Input_Signal,
       ins(14) => Dangling_Input_Signal,
       ins(15) => Dangling_Input_Signal,
       ins(16) => Dangling_Input_Signal,
       ins(17) => Dangling_Input_Signal,
       ins(18) => Dangling_Input_Signal,
       ins(19) => Dangling_Input_Signal,
       ins(20) => Dangling_Input_Signal,
       ins(21) => Dangling_Input_Signal,
       ins(22) => Dangling_Input_Signal,
       ins(23) => Dangling_Input_Signal,
       ins(24) => NET180,
       old_ins(0) => Dangling_Input_Signal,
       old_ins(1) => Dangling_Input_Signal,
       old_ins(2) => Dangling_Input_Signal,
       old_ins(3) => Dangling_Input_Signal,
       old_ins(4) => Dangling_Input_Signal,
       old_ins(5) => Dangling_Input_Signal,
       old_ins(6) => Dangling_Input_Signal,
       old_ins(7) => Dangling_Input_Signal,
       old_ins(8) => Dangling_Input_Signal,
       old_ins(9) => Dangling_Input_Signal,
       old_ins(10) => Dangling_Input_Signal,
       old_ins(11) => Dangling_Input_Signal,
       old_ins(12) => Dangling_Input_Signal,
       old_ins(13) => Dangling_Input_Signal,
       old_ins(14) => Dangling_Input_Signal,
       old_ins(15) => Dangling_Input_Signal,
       old_ins(16) => Dangling_Input_Signal,
       old_ins(17) => Dangling_Input_Signal,
       old_ins(18) => Dangling_Input_Signal,
       old_ins(19) => Dangling_Input_Signal,
       old_ins(20) => Dangling_Input_Signal,
       old_ins(21) => Dangling_Input_Signal,
       old_ins(22) => Dangling_Input_Signal,
       old_ins(23) => Dangling_Input_Signal,
       old_ins(24) => NET246,
       r1_in(0) => Dangling_Input_Signal,
       r1_in(1) => Dangling_Input_Signal,
       r1_in(2) => Dangling_Input_Signal,
       r1_in(3) => Dangling_Input_Signal,
       r1_in(4) => Dangling_Input_Signal,
       r1_in(5) => Dangling_Input_Signal,
       r1_in(6) => Dangling_Input_Signal,
       r1_in(7) => Dangling_Input_Signal,
       r1_in(8) => Dangling_Input_Signal,
       r1_in(9) => Dangling_Input_Signal,
       r1_in(10) => Dangling_Input_Signal,
       r1_in(11) => Dangling_Input_Signal,
       r1_in(12) => Dangling_Input_Signal,
       r1_in(13) => Dangling_Input_Signal,
       r1_in(14) => Dangling_Input_Signal,
       r1_in(15) => Dangling_Input_Signal,
       r1_in(16) => Dangling_Input_Signal,
       r1_in(17) => Dangling_Input_Signal,
       r1_in(18) => Dangling_Input_Signal,
       r1_in(19) => Dangling_Input_Signal,
       r1_in(20) => Dangling_Input_Signal,
       r1_in(21) => Dangling_Input_Signal,
       r1_in(22) => Dangling_Input_Signal,
       r1_in(23) => Dangling_Input_Signal,
       r1_in(24) => Dangling_Input_Signal,
       r1_in(25) => Dangling_Input_Signal,
       r1_in(26) => Dangling_Input_Signal,
       r1_in(27) => Dangling_Input_Signal,
       r1_in(28) => Dangling_Input_Signal,
       r1_in(29) => Dangling_Input_Signal,
       r1_in(30) => Dangling_Input_Signal,
       r1_in(31) => Dangling_Input_Signal,
       r1_in(32) => Dangling_Input_Signal,
       r1_in(33) => Dangling_Input_Signal,
       r1_in(34) => Dangling_Input_Signal,
       r1_in(35) => Dangling_Input_Signal,
       r1_in(36) => Dangling_Input_Signal,
       r1_in(37) => Dangling_Input_Signal,
       r1_in(38) => Dangling_Input_Signal,
       r1_in(39) => Dangling_Input_Signal,
       r1_in(40) => Dangling_Input_Signal,
       r1_in(41) => Dangling_Input_Signal,
       r1_in(42) => Dangling_Input_Signal,
       r1_in(43) => Dangling_Input_Signal,
       r1_in(44) => Dangling_Input_Signal,
       r1_in(45) => Dangling_Input_Signal,
       r1_in(46) => Dangling_Input_Signal,
       r1_in(47) => Dangling_Input_Signal,
       r1_in(48) => Dangling_Input_Signal,
       r1_in(49) => Dangling_Input_Signal,
       r1_in(50) => Dangling_Input_Signal,
       r1_in(51) => Dangling_Input_Signal,
       r1_in(52) => Dangling_Input_Signal,
       r1_in(53) => Dangling_Input_Signal,
       r1_in(54) => Dangling_Input_Signal,
       r1_in(55) => Dangling_Input_Signal,
       r1_in(56) => Dangling_Input_Signal,
       r1_in(57) => Dangling_Input_Signal,
       r1_in(58) => Dangling_Input_Signal,
       r1_in(59) => Dangling_Input_Signal,
       r1_in(60) => Dangling_Input_Signal,
       r1_in(61) => Dangling_Input_Signal,
       r1_in(62) => Dangling_Input_Signal,
       r1_in(63) => Dangling_Input_Signal,
       r1_in(64) => Dangling_Input_Signal,
       r1_in(65) => Dangling_Input_Signal,
       r1_in(66) => Dangling_Input_Signal,
       r1_in(67) => Dangling_Input_Signal,
       r1_in(68) => Dangling_Input_Signal,
       r1_in(69) => Dangling_Input_Signal,
       r1_in(70) => Dangling_Input_Signal,
       r1_in(71) => Dangling_Input_Signal,
       r1_in(72) => Dangling_Input_Signal,
       r1_in(73) => Dangling_Input_Signal,
       r1_in(74) => Dangling_Input_Signal,
       r1_in(75) => Dangling_Input_Signal,
       r1_in(76) => Dangling_Input_Signal,
       r1_in(77) => Dangling_Input_Signal,
       r1_in(78) => Dangling_Input_Signal,
       r1_in(79) => Dangling_Input_Signal,
       r1_in(80) => Dangling_Input_Signal,
       r1_in(81) => Dangling_Input_Signal,
       r1_in(82) => Dangling_Input_Signal,
       r1_in(83) => Dangling_Input_Signal,
       r1_in(84) => Dangling_Input_Signal,
       r1_in(85) => Dangling_Input_Signal,
       r1_in(86) => Dangling_Input_Signal,
       r1_in(87) => Dangling_Input_Signal,
       r1_in(88) => Dangling_Input_Signal,
       r1_in(89) => Dangling_Input_Signal,
       r1_in(90) => Dangling_Input_Signal,
       r1_in(91) => Dangling_Input_Signal,
       r1_in(92) => Dangling_Input_Signal,
       r1_in(93) => Dangling_Input_Signal,
       r1_in(94) => Dangling_Input_Signal,
       r1_in(95) => Dangling_Input_Signal,
       r1_in(96) => Dangling_Input_Signal,
       r1_in(97) => Dangling_Input_Signal,
       r1_in(98) => Dangling_Input_Signal,
       r1_in(99) => Dangling_Input_Signal,
       r1_in(100) => Dangling_Input_Signal,
       r1_in(101) => Dangling_Input_Signal,
       r1_in(102) => Dangling_Input_Signal,
       r1_in(103) => Dangling_Input_Signal,
       r1_in(104) => Dangling_Input_Signal,
       r1_in(105) => Dangling_Input_Signal,
       r1_in(106) => Dangling_Input_Signal,
       r1_in(107) => Dangling_Input_Signal,
       r1_in(108) => Dangling_Input_Signal,
       r1_in(109) => Dangling_Input_Signal,
       r1_in(110) => Dangling_Input_Signal,
       r1_in(111) => Dangling_Input_Signal,
       r1_in(112) => Dangling_Input_Signal,
       r1_in(113) => Dangling_Input_Signal,
       r1_in(114) => Dangling_Input_Signal,
       r1_in(115) => Dangling_Input_Signal,
       r1_in(116) => Dangling_Input_Signal,
       r1_in(117) => Dangling_Input_Signal,
       r1_in(118) => Dangling_Input_Signal,
       r1_in(119) => Dangling_Input_Signal,
       r1_in(120) => Dangling_Input_Signal,
       r1_in(121) => Dangling_Input_Signal,
       r1_in(122) => Dangling_Input_Signal,
       r1_in(123) => Dangling_Input_Signal,
       r1_in(124) => Dangling_Input_Signal,
       r1_in(125) => Dangling_Input_Signal,
       r1_in(126) => Dangling_Input_Signal,
       r1_in(127) => NET122,
       r1_out(0) => DANGLING_U3_r1_out_0,
       r1_out(1) => DANGLING_U3_r1_out_1,
       r1_out(2) => DANGLING_U3_r1_out_2,
       r1_out(3) => DANGLING_U3_r1_out_3,
       r1_out(4) => DANGLING_U3_r1_out_4,
       r1_out(5) => DANGLING_U3_r1_out_5,
       r1_out(6) => DANGLING_U3_r1_out_6,
       r1_out(7) => DANGLING_U3_r1_out_7,
       r1_out(8) => DANGLING_U3_r1_out_8,
       r1_out(9) => DANGLING_U3_r1_out_9,
       r1_out(10) => DANGLING_U3_r1_out_10,
       r1_out(11) => DANGLING_U3_r1_out_11,
       r1_out(12) => DANGLING_U3_r1_out_12,
       r1_out(13) => DANGLING_U3_r1_out_13,
       r1_out(14) => DANGLING_U3_r1_out_14,
       r1_out(15) => DANGLING_U3_r1_out_15,
       r1_out(16) => DANGLING_U3_r1_out_16,
       r1_out(17) => DANGLING_U3_r1_out_17,
       r1_out(18) => DANGLING_U3_r1_out_18,
       r1_out(19) => DANGLING_U3_r1_out_19,
       r1_out(20) => DANGLING_U3_r1_out_20,
       r1_out(21) => DANGLING_U3_r1_out_21,
       r1_out(22) => DANGLING_U3_r1_out_22,
       r1_out(23) => DANGLING_U3_r1_out_23,
       r1_out(24) => DANGLING_U3_r1_out_24,
       r1_out(25) => DANGLING_U3_r1_out_25,
       r1_out(26) => DANGLING_U3_r1_out_26,
       r1_out(27) => DANGLING_U3_r1_out_27,
       r1_out(28) => DANGLING_U3_r1_out_28,
       r1_out(29) => DANGLING_U3_r1_out_29,
       r1_out(30) => DANGLING_U3_r1_out_30,
       r1_out(31) => DANGLING_U3_r1_out_31,
       r1_out(32) => DANGLING_U3_r1_out_32,
       r1_out(33) => DANGLING_U3_r1_out_33,
       r1_out(34) => DANGLING_U3_r1_out_34,
       r1_out(35) => DANGLING_U3_r1_out_35,
       r1_out(36) => DANGLING_U3_r1_out_36,
       r1_out(37) => DANGLING_U3_r1_out_37,
       r1_out(38) => DANGLING_U3_r1_out_38,
       r1_out(39) => DANGLING_U3_r1_out_39,
       r1_out(40) => DANGLING_U3_r1_out_40,
       r1_out(41) => DANGLING_U3_r1_out_41,
       r1_out(42) => DANGLING_U3_r1_out_42,
       r1_out(43) => DANGLING_U3_r1_out_43,
       r1_out(44) => DANGLING_U3_r1_out_44,
       r1_out(45) => DANGLING_U3_r1_out_45,
       r1_out(46) => DANGLING_U3_r1_out_46,
       r1_out(47) => DANGLING_U3_r1_out_47,
       r1_out(48) => DANGLING_U3_r1_out_48,
       r1_out(49) => DANGLING_U3_r1_out_49,
       r1_out(50) => DANGLING_U3_r1_out_50,
       r1_out(51) => DANGLING_U3_r1_out_51,
       r1_out(52) => DANGLING_U3_r1_out_52,
       r1_out(53) => DANGLING_U3_r1_out_53,
       r1_out(54) => DANGLING_U3_r1_out_54,
       r1_out(55) => DANGLING_U3_r1_out_55,
       r1_out(56) => DANGLING_U3_r1_out_56,
       r1_out(57) => DANGLING_U3_r1_out_57,
       r1_out(58) => DANGLING_U3_r1_out_58,
       r1_out(59) => DANGLING_U3_r1_out_59,
       r1_out(60) => DANGLING_U3_r1_out_60,
       r1_out(61) => DANGLING_U3_r1_out_61,
       r1_out(62) => DANGLING_U3_r1_out_62,
       r1_out(63) => DANGLING_U3_r1_out_63,
       r1_out(64) => DANGLING_U3_r1_out_64,
       r1_out(65) => DANGLING_U3_r1_out_65,
       r1_out(66) => DANGLING_U3_r1_out_66,
       r1_out(67) => DANGLING_U3_r1_out_67,
       r1_out(68) => DANGLING_U3_r1_out_68,
       r1_out(69) => DANGLING_U3_r1_out_69,
       r1_out(70) => DANGLING_U3_r1_out_70,
       r1_out(71) => DANGLING_U3_r1_out_71,
       r1_out(72) => DANGLING_U3_r1_out_72,
       r1_out(73) => DANGLING_U3_r1_out_73,
       r1_out(74) => DANGLING_U3_r1_out_74,
       r1_out(75) => DANGLING_U3_r1_out_75,
       r1_out(76) => DANGLING_U3_r1_out_76,
       r1_out(77) => DANGLING_U3_r1_out_77,
       r1_out(78) => DANGLING_U3_r1_out_78,
       r1_out(79) => DANGLING_U3_r1_out_79,
       r1_out(80) => DANGLING_U3_r1_out_80,
       r1_out(81) => DANGLING_U3_r1_out_81,
       r1_out(82) => DANGLING_U3_r1_out_82,
       r1_out(83) => DANGLING_U3_r1_out_83,
       r1_out(84) => DANGLING_U3_r1_out_84,
       r1_out(85) => DANGLING_U3_r1_out_85,
       r1_out(86) => DANGLING_U3_r1_out_86,
       r1_out(87) => DANGLING_U3_r1_out_87,
       r1_out(88) => DANGLING_U3_r1_out_88,
       r1_out(89) => DANGLING_U3_r1_out_89,
       r1_out(90) => DANGLING_U3_r1_out_90,
       r1_out(91) => DANGLING_U3_r1_out_91,
       r1_out(92) => DANGLING_U3_r1_out_92,
       r1_out(93) => DANGLING_U3_r1_out_93,
       r1_out(94) => DANGLING_U3_r1_out_94,
       r1_out(95) => DANGLING_U3_r1_out_95,
       r1_out(96) => DANGLING_U3_r1_out_96,
       r1_out(97) => DANGLING_U3_r1_out_97,
       r1_out(98) => DANGLING_U3_r1_out_98,
       r1_out(99) => DANGLING_U3_r1_out_99,
       r1_out(100) => DANGLING_U3_r1_out_100,
       r1_out(101) => DANGLING_U3_r1_out_101,
       r1_out(102) => DANGLING_U3_r1_out_102,
       r1_out(103) => DANGLING_U3_r1_out_103,
       r1_out(104) => DANGLING_U3_r1_out_104,
       r1_out(105) => DANGLING_U3_r1_out_105,
       r1_out(106) => DANGLING_U3_r1_out_106,
       r1_out(107) => DANGLING_U3_r1_out_107,
       r1_out(108) => DANGLING_U3_r1_out_108,
       r1_out(109) => DANGLING_U3_r1_out_109,
       r1_out(110) => DANGLING_U3_r1_out_110,
       r1_out(111) => DANGLING_U3_r1_out_111,
       r1_out(112) => DANGLING_U3_r1_out_112,
       r1_out(113) => DANGLING_U3_r1_out_113,
       r1_out(114) => DANGLING_U3_r1_out_114,
       r1_out(115) => DANGLING_U3_r1_out_115,
       r1_out(116) => DANGLING_U3_r1_out_116,
       r1_out(117) => DANGLING_U3_r1_out_117,
       r1_out(118) => DANGLING_U3_r1_out_118,
       r1_out(119) => DANGLING_U3_r1_out_119,
       r1_out(120) => DANGLING_U3_r1_out_120,
       r1_out(121) => DANGLING_U3_r1_out_121,
       r1_out(122) => DANGLING_U3_r1_out_122,
       r1_out(123) => DANGLING_U3_r1_out_123,
       r1_out(124) => DANGLING_U3_r1_out_124,
       r1_out(125) => DANGLING_U3_r1_out_125,
       r1_out(126) => DANGLING_U3_r1_out_126,
       r1_out(127) => NET238,
       r2_in(0) => Dangling_Input_Signal,
       r2_in(1) => Dangling_Input_Signal,
       r2_in(2) => Dangling_Input_Signal,
       r2_in(3) => Dangling_Input_Signal,
       r2_in(4) => Dangling_Input_Signal,
       r2_in(5) => Dangling_Input_Signal,
       r2_in(6) => Dangling_Input_Signal,
       r2_in(7) => Dangling_Input_Signal,
       r2_in(8) => Dangling_Input_Signal,
       r2_in(9) => Dangling_Input_Signal,
       r2_in(10) => Dangling_Input_Signal,
       r2_in(11) => Dangling_Input_Signal,
       r2_in(12) => Dangling_Input_Signal,
       r2_in(13) => Dangling_Input_Signal,
       r2_in(14) => Dangling_Input_Signal,
       r2_in(15) => Dangling_Input_Signal,
       r2_in(16) => Dangling_Input_Signal,
       r2_in(17) => Dangling_Input_Signal,
       r2_in(18) => Dangling_Input_Signal,
       r2_in(19) => Dangling_Input_Signal,
       r2_in(20) => Dangling_Input_Signal,
       r2_in(21) => Dangling_Input_Signal,
       r2_in(22) => Dangling_Input_Signal,
       r2_in(23) => Dangling_Input_Signal,
       r2_in(24) => Dangling_Input_Signal,
       r2_in(25) => Dangling_Input_Signal,
       r2_in(26) => Dangling_Input_Signal,
       r2_in(27) => Dangling_Input_Signal,
       r2_in(28) => Dangling_Input_Signal,
       r2_in(29) => Dangling_Input_Signal,
       r2_in(30) => Dangling_Input_Signal,
       r2_in(31) => Dangling_Input_Signal,
       r2_in(32) => Dangling_Input_Signal,
       r2_in(33) => Dangling_Input_Signal,
       r2_in(34) => Dangling_Input_Signal,
       r2_in(35) => Dangling_Input_Signal,
       r2_in(36) => Dangling_Input_Signal,
       r2_in(37) => Dangling_Input_Signal,
       r2_in(38) => Dangling_Input_Signal,
       r2_in(39) => Dangling_Input_Signal,
       r2_in(40) => Dangling_Input_Signal,
       r2_in(41) => Dangling_Input_Signal,
       r2_in(42) => Dangling_Input_Signal,
       r2_in(43) => Dangling_Input_Signal,
       r2_in(44) => Dangling_Input_Signal,
       r2_in(45) => Dangling_Input_Signal,
       r2_in(46) => Dangling_Input_Signal,
       r2_in(47) => Dangling_Input_Signal,
       r2_in(48) => Dangling_Input_Signal,
       r2_in(49) => Dangling_Input_Signal,
       r2_in(50) => Dangling_Input_Signal,
       r2_in(51) => Dangling_Input_Signal,
       r2_in(52) => Dangling_Input_Signal,
       r2_in(53) => Dangling_Input_Signal,
       r2_in(54) => Dangling_Input_Signal,
       r2_in(55) => Dangling_Input_Signal,
       r2_in(56) => Dangling_Input_Signal,
       r2_in(57) => Dangling_Input_Signal,
       r2_in(58) => Dangling_Input_Signal,
       r2_in(59) => Dangling_Input_Signal,
       r2_in(60) => Dangling_Input_Signal,
       r2_in(61) => Dangling_Input_Signal,
       r2_in(62) => Dangling_Input_Signal,
       r2_in(63) => Dangling_Input_Signal,
       r2_in(64) => Dangling_Input_Signal,
       r2_in(65) => Dangling_Input_Signal,
       r2_in(66) => Dangling_Input_Signal,
       r2_in(67) => Dangling_Input_Signal,
       r2_in(68) => Dangling_Input_Signal,
       r2_in(69) => Dangling_Input_Signal,
       r2_in(70) => Dangling_Input_Signal,
       r2_in(71) => Dangling_Input_Signal,
       r2_in(72) => Dangling_Input_Signal,
       r2_in(73) => Dangling_Input_Signal,
       r2_in(74) => Dangling_Input_Signal,
       r2_in(75) => Dangling_Input_Signal,
       r2_in(76) => Dangling_Input_Signal,
       r2_in(77) => Dangling_Input_Signal,
       r2_in(78) => Dangling_Input_Signal,
       r2_in(79) => Dangling_Input_Signal,
       r2_in(80) => Dangling_Input_Signal,
       r2_in(81) => Dangling_Input_Signal,
       r2_in(82) => Dangling_Input_Signal,
       r2_in(83) => Dangling_Input_Signal,
       r2_in(84) => Dangling_Input_Signal,
       r2_in(85) => Dangling_Input_Signal,
       r2_in(86) => Dangling_Input_Signal,
       r2_in(87) => Dangling_Input_Signal,
       r2_in(88) => Dangling_Input_Signal,
       r2_in(89) => Dangling_Input_Signal,
       r2_in(90) => Dangling_Input_Signal,
       r2_in(91) => Dangling_Input_Signal,
       r2_in(92) => Dangling_Input_Signal,
       r2_in(93) => Dangling_Input_Signal,
       r2_in(94) => Dangling_Input_Signal,
       r2_in(95) => Dangling_Input_Signal,
       r2_in(96) => Dangling_Input_Signal,
       r2_in(97) => Dangling_Input_Signal,
       r2_in(98) => Dangling_Input_Signal,
       r2_in(99) => Dangling_Input_Signal,
       r2_in(100) => Dangling_Input_Signal,
       r2_in(101) => Dangling_Input_Signal,
       r2_in(102) => Dangling_Input_Signal,
       r2_in(103) => Dangling_Input_Signal,
       r2_in(104) => Dangling_Input_Signal,
       r2_in(105) => Dangling_Input_Signal,
       r2_in(106) => Dangling_Input_Signal,
       r2_in(107) => Dangling_Input_Signal,
       r2_in(108) => Dangling_Input_Signal,
       r2_in(109) => Dangling_Input_Signal,
       r2_in(110) => Dangling_Input_Signal,
       r2_in(111) => Dangling_Input_Signal,
       r2_in(112) => Dangling_Input_Signal,
       r2_in(113) => Dangling_Input_Signal,
       r2_in(114) => Dangling_Input_Signal,
       r2_in(115) => Dangling_Input_Signal,
       r2_in(116) => Dangling_Input_Signal,
       r2_in(117) => Dangling_Input_Signal,
       r2_in(118) => Dangling_Input_Signal,
       r2_in(119) => Dangling_Input_Signal,
       r2_in(120) => Dangling_Input_Signal,
       r2_in(121) => Dangling_Input_Signal,
       r2_in(122) => Dangling_Input_Signal,
       r2_in(123) => Dangling_Input_Signal,
       r2_in(124) => Dangling_Input_Signal,
       r2_in(125) => Dangling_Input_Signal,
       r2_in(126) => Dangling_Input_Signal,
       r2_in(127) => NET134,
       r2_out(0) => DANGLING_U3_r2_out_0,
       r2_out(1) => DANGLING_U3_r2_out_1,
       r2_out(2) => DANGLING_U3_r2_out_2,
       r2_out(3) => DANGLING_U3_r2_out_3,
       r2_out(4) => DANGLING_U3_r2_out_4,
       r2_out(5) => DANGLING_U3_r2_out_5,
       r2_out(6) => DANGLING_U3_r2_out_6,
       r2_out(7) => DANGLING_U3_r2_out_7,
       r2_out(8) => DANGLING_U3_r2_out_8,
       r2_out(9) => DANGLING_U3_r2_out_9,
       r2_out(10) => DANGLING_U3_r2_out_10,
       r2_out(11) => DANGLING_U3_r2_out_11,
       r2_out(12) => DANGLING_U3_r2_out_12,
       r2_out(13) => DANGLING_U3_r2_out_13,
       r2_out(14) => DANGLING_U3_r2_out_14,
       r2_out(15) => DANGLING_U3_r2_out_15,
       r2_out(16) => DANGLING_U3_r2_out_16,
       r2_out(17) => DANGLING_U3_r2_out_17,
       r2_out(18) => DANGLING_U3_r2_out_18,
       r2_out(19) => DANGLING_U3_r2_out_19,
       r2_out(20) => DANGLING_U3_r2_out_20,
       r2_out(21) => DANGLING_U3_r2_out_21,
       r2_out(22) => DANGLING_U3_r2_out_22,
       r2_out(23) => DANGLING_U3_r2_out_23,
       r2_out(24) => DANGLING_U3_r2_out_24,
       r2_out(25) => DANGLING_U3_r2_out_25,
       r2_out(26) => DANGLING_U3_r2_out_26,
       r2_out(27) => DANGLING_U3_r2_out_27,
       r2_out(28) => DANGLING_U3_r2_out_28,
       r2_out(29) => DANGLING_U3_r2_out_29,
       r2_out(30) => DANGLING_U3_r2_out_30,
       r2_out(31) => DANGLING_U3_r2_out_31,
       r2_out(32) => DANGLING_U3_r2_out_32,
       r2_out(33) => DANGLING_U3_r2_out_33,
       r2_out(34) => DANGLING_U3_r2_out_34,
       r2_out(35) => DANGLING_U3_r2_out_35,
       r2_out(36) => DANGLING_U3_r2_out_36,
       r2_out(37) => DANGLING_U3_r2_out_37,
       r2_out(38) => DANGLING_U3_r2_out_38,
       r2_out(39) => DANGLING_U3_r2_out_39,
       r2_out(40) => DANGLING_U3_r2_out_40,
       r2_out(41) => DANGLING_U3_r2_out_41,
       r2_out(42) => DANGLING_U3_r2_out_42,
       r2_out(43) => DANGLING_U3_r2_out_43,
       r2_out(44) => DANGLING_U3_r2_out_44,
       r2_out(45) => DANGLING_U3_r2_out_45,
       r2_out(46) => DANGLING_U3_r2_out_46,
       r2_out(47) => DANGLING_U3_r2_out_47,
       r2_out(48) => DANGLING_U3_r2_out_48,
       r2_out(49) => DANGLING_U3_r2_out_49,
       r2_out(50) => DANGLING_U3_r2_out_50,
       r2_out(51) => DANGLING_U3_r2_out_51,
       r2_out(52) => DANGLING_U3_r2_out_52,
       r2_out(53) => DANGLING_U3_r2_out_53,
       r2_out(54) => DANGLING_U3_r2_out_54,
       r2_out(55) => DANGLING_U3_r2_out_55,
       r2_out(56) => DANGLING_U3_r2_out_56,
       r2_out(57) => DANGLING_U3_r2_out_57,
       r2_out(58) => DANGLING_U3_r2_out_58,
       r2_out(59) => DANGLING_U3_r2_out_59,
       r2_out(60) => DANGLING_U3_r2_out_60,
       r2_out(61) => DANGLING_U3_r2_out_61,
       r2_out(62) => DANGLING_U3_r2_out_62,
       r2_out(63) => DANGLING_U3_r2_out_63,
       r2_out(64) => DANGLING_U3_r2_out_64,
       r2_out(65) => DANGLING_U3_r2_out_65,
       r2_out(66) => DANGLING_U3_r2_out_66,
       r2_out(67) => DANGLING_U3_r2_out_67,
       r2_out(68) => DANGLING_U3_r2_out_68,
       r2_out(69) => DANGLING_U3_r2_out_69,
       r2_out(70) => DANGLING_U3_r2_out_70,
       r2_out(71) => DANGLING_U3_r2_out_71,
       r2_out(72) => DANGLING_U3_r2_out_72,
       r2_out(73) => DANGLING_U3_r2_out_73,
       r2_out(74) => DANGLING_U3_r2_out_74,
       r2_out(75) => DANGLING_U3_r2_out_75,
       r2_out(76) => DANGLING_U3_r2_out_76,
       r2_out(77) => DANGLING_U3_r2_out_77,
       r2_out(78) => DANGLING_U3_r2_out_78,
       r2_out(79) => DANGLING_U3_r2_out_79,
       r2_out(80) => DANGLING_U3_r2_out_80,
       r2_out(81) => DANGLING_U3_r2_out_81,
       r2_out(82) => DANGLING_U3_r2_out_82,
       r2_out(83) => DANGLING_U3_r2_out_83,
       r2_out(84) => DANGLING_U3_r2_out_84,
       r2_out(85) => DANGLING_U3_r2_out_85,
       r2_out(86) => DANGLING_U3_r2_out_86,
       r2_out(87) => DANGLING_U3_r2_out_87,
       r2_out(88) => DANGLING_U3_r2_out_88,
       r2_out(89) => DANGLING_U3_r2_out_89,
       r2_out(90) => DANGLING_U3_r2_out_90,
       r2_out(91) => DANGLING_U3_r2_out_91,
       r2_out(92) => DANGLING_U3_r2_out_92,
       r2_out(93) => DANGLING_U3_r2_out_93,
       r2_out(94) => DANGLING_U3_r2_out_94,
       r2_out(95) => DANGLING_U3_r2_out_95,
       r2_out(96) => DANGLING_U3_r2_out_96,
       r2_out(97) => DANGLING_U3_r2_out_97,
       r2_out(98) => DANGLING_U3_r2_out_98,
       r2_out(99) => DANGLING_U3_r2_out_99,
       r2_out(100) => DANGLING_U3_r2_out_100,
       r2_out(101) => DANGLING_U3_r2_out_101,
       r2_out(102) => DANGLING_U3_r2_out_102,
       r2_out(103) => DANGLING_U3_r2_out_103,
       r2_out(104) => DANGLING_U3_r2_out_104,
       r2_out(105) => DANGLING_U3_r2_out_105,
       r2_out(106) => DANGLING_U3_r2_out_106,
       r2_out(107) => DANGLING_U3_r2_out_107,
       r2_out(108) => DANGLING_U3_r2_out_108,
       r2_out(109) => DANGLING_U3_r2_out_109,
       r2_out(110) => DANGLING_U3_r2_out_110,
       r2_out(111) => DANGLING_U3_r2_out_111,
       r2_out(112) => DANGLING_U3_r2_out_112,
       r2_out(113) => DANGLING_U3_r2_out_113,
       r2_out(114) => DANGLING_U3_r2_out_114,
       r2_out(115) => DANGLING_U3_r2_out_115,
       r2_out(116) => DANGLING_U3_r2_out_116,
       r2_out(117) => DANGLING_U3_r2_out_117,
       r2_out(118) => DANGLING_U3_r2_out_118,
       r2_out(119) => DANGLING_U3_r2_out_119,
       r2_out(120) => DANGLING_U3_r2_out_120,
       r2_out(121) => DANGLING_U3_r2_out_121,
       r2_out(122) => DANGLING_U3_r2_out_122,
       r2_out(123) => DANGLING_U3_r2_out_123,
       r2_out(124) => DANGLING_U3_r2_out_124,
       r2_out(125) => DANGLING_U3_r2_out_125,
       r2_out(126) => DANGLING_U3_r2_out_126,
       r2_out(127) => NET230,
       r3_in(0) => Dangling_Input_Signal,
       r3_in(1) => Dangling_Input_Signal,
       r3_in(2) => Dangling_Input_Signal,
       r3_in(3) => Dangling_Input_Signal,
       r3_in(4) => Dangling_Input_Signal,
       r3_in(5) => Dangling_Input_Signal,
       r3_in(6) => Dangling_Input_Signal,
       r3_in(7) => Dangling_Input_Signal,
       r3_in(8) => Dangling_Input_Signal,
       r3_in(9) => Dangling_Input_Signal,
       r3_in(10) => Dangling_Input_Signal,
       r3_in(11) => Dangling_Input_Signal,
       r3_in(12) => Dangling_Input_Signal,
       r3_in(13) => Dangling_Input_Signal,
       r3_in(14) => Dangling_Input_Signal,
       r3_in(15) => Dangling_Input_Signal,
       r3_in(16) => Dangling_Input_Signal,
       r3_in(17) => Dangling_Input_Signal,
       r3_in(18) => Dangling_Input_Signal,
       r3_in(19) => Dangling_Input_Signal,
       r3_in(20) => Dangling_Input_Signal,
       r3_in(21) => Dangling_Input_Signal,
       r3_in(22) => Dangling_Input_Signal,
       r3_in(23) => Dangling_Input_Signal,
       r3_in(24) => Dangling_Input_Signal,
       r3_in(25) => Dangling_Input_Signal,
       r3_in(26) => Dangling_Input_Signal,
       r3_in(27) => Dangling_Input_Signal,
       r3_in(28) => Dangling_Input_Signal,
       r3_in(29) => Dangling_Input_Signal,
       r3_in(30) => Dangling_Input_Signal,
       r3_in(31) => Dangling_Input_Signal,
       r3_in(32) => Dangling_Input_Signal,
       r3_in(33) => Dangling_Input_Signal,
       r3_in(34) => Dangling_Input_Signal,
       r3_in(35) => Dangling_Input_Signal,
       r3_in(36) => Dangling_Input_Signal,
       r3_in(37) => Dangling_Input_Signal,
       r3_in(38) => Dangling_Input_Signal,
       r3_in(39) => Dangling_Input_Signal,
       r3_in(40) => Dangling_Input_Signal,
       r3_in(41) => Dangling_Input_Signal,
       r3_in(42) => Dangling_Input_Signal,
       r3_in(43) => Dangling_Input_Signal,
       r3_in(44) => Dangling_Input_Signal,
       r3_in(45) => Dangling_Input_Signal,
       r3_in(46) => Dangling_Input_Signal,
       r3_in(47) => Dangling_Input_Signal,
       r3_in(48) => Dangling_Input_Signal,
       r3_in(49) => Dangling_Input_Signal,
       r3_in(50) => Dangling_Input_Signal,
       r3_in(51) => Dangling_Input_Signal,
       r3_in(52) => Dangling_Input_Signal,
       r3_in(53) => Dangling_Input_Signal,
       r3_in(54) => Dangling_Input_Signal,
       r3_in(55) => Dangling_Input_Signal,
       r3_in(56) => Dangling_Input_Signal,
       r3_in(57) => Dangling_Input_Signal,
       r3_in(58) => Dangling_Input_Signal,
       r3_in(59) => Dangling_Input_Signal,
       r3_in(60) => Dangling_Input_Signal,
       r3_in(61) => Dangling_Input_Signal,
       r3_in(62) => Dangling_Input_Signal,
       r3_in(63) => Dangling_Input_Signal,
       r3_in(64) => Dangling_Input_Signal,
       r3_in(65) => Dangling_Input_Signal,
       r3_in(66) => Dangling_Input_Signal,
       r3_in(67) => Dangling_Input_Signal,
       r3_in(68) => Dangling_Input_Signal,
       r3_in(69) => Dangling_Input_Signal,
       r3_in(70) => Dangling_Input_Signal,
       r3_in(71) => Dangling_Input_Signal,
       r3_in(72) => Dangling_Input_Signal,
       r3_in(73) => Dangling_Input_Signal,
       r3_in(74) => Dangling_Input_Signal,
       r3_in(75) => Dangling_Input_Signal,
       r3_in(76) => Dangling_Input_Signal,
       r3_in(77) => Dangling_Input_Signal,
       r3_in(78) => Dangling_Input_Signal,
       r3_in(79) => Dangling_Input_Signal,
       r3_in(80) => Dangling_Input_Signal,
       r3_in(81) => Dangling_Input_Signal,
       r3_in(82) => Dangling_Input_Signal,
       r3_in(83) => Dangling_Input_Signal,
       r3_in(84) => Dangling_Input_Signal,
       r3_in(85) => Dangling_Input_Signal,
       r3_in(86) => Dangling_Input_Signal,
       r3_in(87) => Dangling_Input_Signal,
       r3_in(88) => Dangling_Input_Signal,
       r3_in(89) => Dangling_Input_Signal,
       r3_in(90) => Dangling_Input_Signal,
       r3_in(91) => Dangling_Input_Signal,
       r3_in(92) => Dangling_Input_Signal,
       r3_in(93) => Dangling_Input_Signal,
       r3_in(94) => Dangling_Input_Signal,
       r3_in(95) => Dangling_Input_Signal,
       r3_in(96) => Dangling_Input_Signal,
       r3_in(97) => Dangling_Input_Signal,
       r3_in(98) => Dangling_Input_Signal,
       r3_in(99) => Dangling_Input_Signal,
       r3_in(100) => Dangling_Input_Signal,
       r3_in(101) => Dangling_Input_Signal,
       r3_in(102) => Dangling_Input_Signal,
       r3_in(103) => Dangling_Input_Signal,
       r3_in(104) => Dangling_Input_Signal,
       r3_in(105) => Dangling_Input_Signal,
       r3_in(106) => Dangling_Input_Signal,
       r3_in(107) => Dangling_Input_Signal,
       r3_in(108) => Dangling_Input_Signal,
       r3_in(109) => Dangling_Input_Signal,
       r3_in(110) => Dangling_Input_Signal,
       r3_in(111) => Dangling_Input_Signal,
       r3_in(112) => Dangling_Input_Signal,
       r3_in(113) => Dangling_Input_Signal,
       r3_in(114) => Dangling_Input_Signal,
       r3_in(115) => Dangling_Input_Signal,
       r3_in(116) => Dangling_Input_Signal,
       r3_in(117) => Dangling_Input_Signal,
       r3_in(118) => Dangling_Input_Signal,
       r3_in(119) => Dangling_Input_Signal,
       r3_in(120) => Dangling_Input_Signal,
       r3_in(121) => Dangling_Input_Signal,
       r3_in(122) => Dangling_Input_Signal,
       r3_in(123) => Dangling_Input_Signal,
       r3_in(124) => Dangling_Input_Signal,
       r3_in(125) => Dangling_Input_Signal,
       r3_in(126) => Dangling_Input_Signal,
       r3_in(127) => NET168,
       r3_out(0) => DANGLING_U3_r3_out_0,
       r3_out(1) => DANGLING_U3_r3_out_1,
       r3_out(2) => DANGLING_U3_r3_out_2,
       r3_out(3) => DANGLING_U3_r3_out_3,
       r3_out(4) => DANGLING_U3_r3_out_4,
       r3_out(5) => DANGLING_U3_r3_out_5,
       r3_out(6) => DANGLING_U3_r3_out_6,
       r3_out(7) => DANGLING_U3_r3_out_7,
       r3_out(8) => DANGLING_U3_r3_out_8,
       r3_out(9) => DANGLING_U3_r3_out_9,
       r3_out(10) => DANGLING_U3_r3_out_10,
       r3_out(11) => DANGLING_U3_r3_out_11,
       r3_out(12) => DANGLING_U3_r3_out_12,
       r3_out(13) => DANGLING_U3_r3_out_13,
       r3_out(14) => DANGLING_U3_r3_out_14,
       r3_out(15) => DANGLING_U3_r3_out_15,
       r3_out(16) => DANGLING_U3_r3_out_16,
       r3_out(17) => DANGLING_U3_r3_out_17,
       r3_out(18) => DANGLING_U3_r3_out_18,
       r3_out(19) => DANGLING_U3_r3_out_19,
       r3_out(20) => DANGLING_U3_r3_out_20,
       r3_out(21) => DANGLING_U3_r3_out_21,
       r3_out(22) => DANGLING_U3_r3_out_22,
       r3_out(23) => DANGLING_U3_r3_out_23,
       r3_out(24) => DANGLING_U3_r3_out_24,
       r3_out(25) => DANGLING_U3_r3_out_25,
       r3_out(26) => DANGLING_U3_r3_out_26,
       r3_out(27) => DANGLING_U3_r3_out_27,
       r3_out(28) => DANGLING_U3_r3_out_28,
       r3_out(29) => DANGLING_U3_r3_out_29,
       r3_out(30) => DANGLING_U3_r3_out_30,
       r3_out(31) => DANGLING_U3_r3_out_31,
       r3_out(32) => DANGLING_U3_r3_out_32,
       r3_out(33) => DANGLING_U3_r3_out_33,
       r3_out(34) => DANGLING_U3_r3_out_34,
       r3_out(35) => DANGLING_U3_r3_out_35,
       r3_out(36) => DANGLING_U3_r3_out_36,
       r3_out(37) => DANGLING_U3_r3_out_37,
       r3_out(38) => DANGLING_U3_r3_out_38,
       r3_out(39) => DANGLING_U3_r3_out_39,
       r3_out(40) => DANGLING_U3_r3_out_40,
       r3_out(41) => DANGLING_U3_r3_out_41,
       r3_out(42) => DANGLING_U3_r3_out_42,
       r3_out(43) => DANGLING_U3_r3_out_43,
       r3_out(44) => DANGLING_U3_r3_out_44,
       r3_out(45) => DANGLING_U3_r3_out_45,
       r3_out(46) => DANGLING_U3_r3_out_46,
       r3_out(47) => DANGLING_U3_r3_out_47,
       r3_out(48) => DANGLING_U3_r3_out_48,
       r3_out(49) => DANGLING_U3_r3_out_49,
       r3_out(50) => DANGLING_U3_r3_out_50,
       r3_out(51) => DANGLING_U3_r3_out_51,
       r3_out(52) => DANGLING_U3_r3_out_52,
       r3_out(53) => DANGLING_U3_r3_out_53,
       r3_out(54) => DANGLING_U3_r3_out_54,
       r3_out(55) => DANGLING_U3_r3_out_55,
       r3_out(56) => DANGLING_U3_r3_out_56,
       r3_out(57) => DANGLING_U3_r3_out_57,
       r3_out(58) => DANGLING_U3_r3_out_58,
       r3_out(59) => DANGLING_U3_r3_out_59,
       r3_out(60) => DANGLING_U3_r3_out_60,
       r3_out(61) => DANGLING_U3_r3_out_61,
       r3_out(62) => DANGLING_U3_r3_out_62,
       r3_out(63) => DANGLING_U3_r3_out_63,
       r3_out(64) => DANGLING_U3_r3_out_64,
       r3_out(65) => DANGLING_U3_r3_out_65,
       r3_out(66) => DANGLING_U3_r3_out_66,
       r3_out(67) => DANGLING_U3_r3_out_67,
       r3_out(68) => DANGLING_U3_r3_out_68,
       r3_out(69) => DANGLING_U3_r3_out_69,
       r3_out(70) => DANGLING_U3_r3_out_70,
       r3_out(71) => DANGLING_U3_r3_out_71,
       r3_out(72) => DANGLING_U3_r3_out_72,
       r3_out(73) => DANGLING_U3_r3_out_73,
       r3_out(74) => DANGLING_U3_r3_out_74,
       r3_out(75) => DANGLING_U3_r3_out_75,
       r3_out(76) => DANGLING_U3_r3_out_76,
       r3_out(77) => DANGLING_U3_r3_out_77,
       r3_out(78) => DANGLING_U3_r3_out_78,
       r3_out(79) => DANGLING_U3_r3_out_79,
       r3_out(80) => DANGLING_U3_r3_out_80,
       r3_out(81) => DANGLING_U3_r3_out_81,
       r3_out(82) => DANGLING_U3_r3_out_82,
       r3_out(83) => DANGLING_U3_r3_out_83,
       r3_out(84) => DANGLING_U3_r3_out_84,
       r3_out(85) => DANGLING_U3_r3_out_85,
       r3_out(86) => DANGLING_U3_r3_out_86,
       r3_out(87) => DANGLING_U3_r3_out_87,
       r3_out(88) => DANGLING_U3_r3_out_88,
       r3_out(89) => DANGLING_U3_r3_out_89,
       r3_out(90) => DANGLING_U3_r3_out_90,
       r3_out(91) => DANGLING_U3_r3_out_91,
       r3_out(92) => DANGLING_U3_r3_out_92,
       r3_out(93) => DANGLING_U3_r3_out_93,
       r3_out(94) => DANGLING_U3_r3_out_94,
       r3_out(95) => DANGLING_U3_r3_out_95,
       r3_out(96) => DANGLING_U3_r3_out_96,
       r3_out(97) => DANGLING_U3_r3_out_97,
       r3_out(98) => DANGLING_U3_r3_out_98,
       r3_out(99) => DANGLING_U3_r3_out_99,
       r3_out(100) => DANGLING_U3_r3_out_100,
       r3_out(101) => DANGLING_U3_r3_out_101,
       r3_out(102) => DANGLING_U3_r3_out_102,
       r3_out(103) => DANGLING_U3_r3_out_103,
       r3_out(104) => DANGLING_U3_r3_out_104,
       r3_out(105) => DANGLING_U3_r3_out_105,
       r3_out(106) => DANGLING_U3_r3_out_106,
       r3_out(107) => DANGLING_U3_r3_out_107,
       r3_out(108) => DANGLING_U3_r3_out_108,
       r3_out(109) => DANGLING_U3_r3_out_109,
       r3_out(110) => DANGLING_U3_r3_out_110,
       r3_out(111) => DANGLING_U3_r3_out_111,
       r3_out(112) => DANGLING_U3_r3_out_112,
       r3_out(113) => DANGLING_U3_r3_out_113,
       r3_out(114) => DANGLING_U3_r3_out_114,
       r3_out(115) => DANGLING_U3_r3_out_115,
       r3_out(116) => DANGLING_U3_r3_out_116,
       r3_out(117) => DANGLING_U3_r3_out_117,
       r3_out(118) => DANGLING_U3_r3_out_118,
       r3_out(119) => DANGLING_U3_r3_out_119,
       r3_out(120) => DANGLING_U3_r3_out_120,
       r3_out(121) => DANGLING_U3_r3_out_121,
       r3_out(122) => DANGLING_U3_r3_out_122,
       r3_out(123) => DANGLING_U3_r3_out_123,
       r3_out(124) => DANGLING_U3_r3_out_124,
       r3_out(125) => DANGLING_U3_r3_out_125,
       r3_out(126) => DANGLING_U3_r3_out_126,
       r3_out(127) => NET222
  );

U5 : register_file
  port map(
       ins(0) => Dangling_Input_Signal,
       ins(1) => Dangling_Input_Signal,
       ins(2) => Dangling_Input_Signal,
       ins(3) => Dangling_Input_Signal,
       ins(4) => Dangling_Input_Signal,
       ins(5) => Dangling_Input_Signal,
       ins(6) => Dangling_Input_Signal,
       ins(7) => Dangling_Input_Signal,
       ins(8) => Dangling_Input_Signal,
       ins(9) => Dangling_Input_Signal,
       ins(10) => Dangling_Input_Signal,
       ins(11) => Dangling_Input_Signal,
       ins(12) => Dangling_Input_Signal,
       ins(13) => Dangling_Input_Signal,
       ins(14) => Dangling_Input_Signal,
       ins(15) => Dangling_Input_Signal,
       ins(16) => Dangling_Input_Signal,
       ins(17) => Dangling_Input_Signal,
       ins(18) => Dangling_Input_Signal,
       ins(19) => Dangling_Input_Signal,
       ins(20) => Dangling_Input_Signal,
       ins(21) => Dangling_Input_Signal,
       ins(22) => Dangling_Input_Signal,
       ins(23) => Dangling_Input_Signal,
       ins(24) => NET114,
       ins_out(0) => DANGLING_U5_ins_out_0,
       ins_out(1) => DANGLING_U5_ins_out_1,
       ins_out(2) => DANGLING_U5_ins_out_2,
       ins_out(3) => DANGLING_U5_ins_out_3,
       ins_out(4) => DANGLING_U5_ins_out_4,
       ins_out(5) => DANGLING_U5_ins_out_5,
       ins_out(6) => DANGLING_U5_ins_out_6,
       ins_out(7) => DANGLING_U5_ins_out_7,
       ins_out(8) => DANGLING_U5_ins_out_8,
       ins_out(9) => DANGLING_U5_ins_out_9,
       ins_out(10) => DANGLING_U5_ins_out_10,
       ins_out(11) => DANGLING_U5_ins_out_11,
       ins_out(12) => DANGLING_U5_ins_out_12,
       ins_out(13) => DANGLING_U5_ins_out_13,
       ins_out(14) => DANGLING_U5_ins_out_14,
       ins_out(15) => DANGLING_U5_ins_out_15,
       ins_out(16) => DANGLING_U5_ins_out_16,
       ins_out(17) => DANGLING_U5_ins_out_17,
       ins_out(18) => DANGLING_U5_ins_out_18,
       ins_out(19) => DANGLING_U5_ins_out_19,
       ins_out(20) => DANGLING_U5_ins_out_20,
       ins_out(21) => DANGLING_U5_ins_out_21,
       ins_out(22) => DANGLING_U5_ins_out_22,
       ins_out(23) => DANGLING_U5_ins_out_23,
       ins_out(24) => NET180,
       old_ins(0) => Dangling_Input_Signal,
       old_ins(1) => Dangling_Input_Signal,
       old_ins(2) => Dangling_Input_Signal,
       old_ins(3) => Dangling_Input_Signal,
       old_ins(4) => Dangling_Input_Signal,
       old_ins(5) => Dangling_Input_Signal,
       old_ins(6) => Dangling_Input_Signal,
       old_ins(7) => Dangling_Input_Signal,
       old_ins(8) => Dangling_Input_Signal,
       old_ins(9) => Dangling_Input_Signal,
       old_ins(10) => Dangling_Input_Signal,
       old_ins(11) => Dangling_Input_Signal,
       old_ins(12) => Dangling_Input_Signal,
       old_ins(13) => Dangling_Input_Signal,
       old_ins(14) => Dangling_Input_Signal,
       old_ins(15) => Dangling_Input_Signal,
       old_ins(16) => Dangling_Input_Signal,
       old_ins(17) => Dangling_Input_Signal,
       old_ins(18) => Dangling_Input_Signal,
       old_ins(19) => Dangling_Input_Signal,
       old_ins(20) => Dangling_Input_Signal,
       old_ins(21) => Dangling_Input_Signal,
       old_ins(22) => Dangling_Input_Signal,
       old_ins(23) => Dangling_Input_Signal,
       old_ins(24) => NET246,
       r1(0) => DANGLING_U5_r1_0,
       r1(1) => DANGLING_U5_r1_1,
       r1(2) => DANGLING_U5_r1_2,
       r1(3) => DANGLING_U5_r1_3,
       r1(4) => DANGLING_U5_r1_4,
       r1(5) => DANGLING_U5_r1_5,
       r1(6) => DANGLING_U5_r1_6,
       r1(7) => DANGLING_U5_r1_7,
       r1(8) => DANGLING_U5_r1_8,
       r1(9) => DANGLING_U5_r1_9,
       r1(10) => DANGLING_U5_r1_10,
       r1(11) => DANGLING_U5_r1_11,
       r1(12) => DANGLING_U5_r1_12,
       r1(13) => DANGLING_U5_r1_13,
       r1(14) => DANGLING_U5_r1_14,
       r1(15) => DANGLING_U5_r1_15,
       r1(16) => DANGLING_U5_r1_16,
       r1(17) => DANGLING_U5_r1_17,
       r1(18) => DANGLING_U5_r1_18,
       r1(19) => DANGLING_U5_r1_19,
       r1(20) => DANGLING_U5_r1_20,
       r1(21) => DANGLING_U5_r1_21,
       r1(22) => DANGLING_U5_r1_22,
       r1(23) => DANGLING_U5_r1_23,
       r1(24) => DANGLING_U5_r1_24,
       r1(25) => DANGLING_U5_r1_25,
       r1(26) => DANGLING_U5_r1_26,
       r1(27) => DANGLING_U5_r1_27,
       r1(28) => DANGLING_U5_r1_28,
       r1(29) => DANGLING_U5_r1_29,
       r1(30) => DANGLING_U5_r1_30,
       r1(31) => DANGLING_U5_r1_31,
       r1(32) => DANGLING_U5_r1_32,
       r1(33) => DANGLING_U5_r1_33,
       r1(34) => DANGLING_U5_r1_34,
       r1(35) => DANGLING_U5_r1_35,
       r1(36) => DANGLING_U5_r1_36,
       r1(37) => DANGLING_U5_r1_37,
       r1(38) => DANGLING_U5_r1_38,
       r1(39) => DANGLING_U5_r1_39,
       r1(40) => DANGLING_U5_r1_40,
       r1(41) => DANGLING_U5_r1_41,
       r1(42) => DANGLING_U5_r1_42,
       r1(43) => DANGLING_U5_r1_43,
       r1(44) => DANGLING_U5_r1_44,
       r1(45) => DANGLING_U5_r1_45,
       r1(46) => DANGLING_U5_r1_46,
       r1(47) => DANGLING_U5_r1_47,
       r1(48) => DANGLING_U5_r1_48,
       r1(49) => DANGLING_U5_r1_49,
       r1(50) => DANGLING_U5_r1_50,
       r1(51) => DANGLING_U5_r1_51,
       r1(52) => DANGLING_U5_r1_52,
       r1(53) => DANGLING_U5_r1_53,
       r1(54) => DANGLING_U5_r1_54,
       r1(55) => DANGLING_U5_r1_55,
       r1(56) => DANGLING_U5_r1_56,
       r1(57) => DANGLING_U5_r1_57,
       r1(58) => DANGLING_U5_r1_58,
       r1(59) => DANGLING_U5_r1_59,
       r1(60) => DANGLING_U5_r1_60,
       r1(61) => DANGLING_U5_r1_61,
       r1(62) => DANGLING_U5_r1_62,
       r1(63) => DANGLING_U5_r1_63,
       r1(64) => DANGLING_U5_r1_64,
       r1(65) => DANGLING_U5_r1_65,
       r1(66) => DANGLING_U5_r1_66,
       r1(67) => DANGLING_U5_r1_67,
       r1(68) => DANGLING_U5_r1_68,
       r1(69) => DANGLING_U5_r1_69,
       r1(70) => DANGLING_U5_r1_70,
       r1(71) => DANGLING_U5_r1_71,
       r1(72) => DANGLING_U5_r1_72,
       r1(73) => DANGLING_U5_r1_73,
       r1(74) => DANGLING_U5_r1_74,
       r1(75) => DANGLING_U5_r1_75,
       r1(76) => DANGLING_U5_r1_76,
       r1(77) => DANGLING_U5_r1_77,
       r1(78) => DANGLING_U5_r1_78,
       r1(79) => DANGLING_U5_r1_79,
       r1(80) => DANGLING_U5_r1_80,
       r1(81) => DANGLING_U5_r1_81,
       r1(82) => DANGLING_U5_r1_82,
       r1(83) => DANGLING_U5_r1_83,
       r1(84) => DANGLING_U5_r1_84,
       r1(85) => DANGLING_U5_r1_85,
       r1(86) => DANGLING_U5_r1_86,
       r1(87) => DANGLING_U5_r1_87,
       r1(88) => DANGLING_U5_r1_88,
       r1(89) => DANGLING_U5_r1_89,
       r1(90) => DANGLING_U5_r1_90,
       r1(91) => DANGLING_U5_r1_91,
       r1(92) => DANGLING_U5_r1_92,
       r1(93) => DANGLING_U5_r1_93,
       r1(94) => DANGLING_U5_r1_94,
       r1(95) => DANGLING_U5_r1_95,
       r1(96) => DANGLING_U5_r1_96,
       r1(97) => DANGLING_U5_r1_97,
       r1(98) => DANGLING_U5_r1_98,
       r1(99) => DANGLING_U5_r1_99,
       r1(100) => DANGLING_U5_r1_100,
       r1(101) => DANGLING_U5_r1_101,
       r1(102) => DANGLING_U5_r1_102,
       r1(103) => DANGLING_U5_r1_103,
       r1(104) => DANGLING_U5_r1_104,
       r1(105) => DANGLING_U5_r1_105,
       r1(106) => DANGLING_U5_r1_106,
       r1(107) => DANGLING_U5_r1_107,
       r1(108) => DANGLING_U5_r1_108,
       r1(109) => DANGLING_U5_r1_109,
       r1(110) => DANGLING_U5_r1_110,
       r1(111) => DANGLING_U5_r1_111,
       r1(112) => DANGLING_U5_r1_112,
       r1(113) => DANGLING_U5_r1_113,
       r1(114) => DANGLING_U5_r1_114,
       r1(115) => DANGLING_U5_r1_115,
       r1(116) => DANGLING_U5_r1_116,
       r1(117) => DANGLING_U5_r1_117,
       r1(118) => DANGLING_U5_r1_118,
       r1(119) => DANGLING_U5_r1_119,
       r1(120) => DANGLING_U5_r1_120,
       r1(121) => DANGLING_U5_r1_121,
       r1(122) => DANGLING_U5_r1_122,
       r1(123) => DANGLING_U5_r1_123,
       r1(124) => DANGLING_U5_r1_124,
       r1(125) => DANGLING_U5_r1_125,
       r1(126) => DANGLING_U5_r1_126,
       r1(127) => NET122,
       r2(0) => DANGLING_U5_r2_0,
       r2(1) => DANGLING_U5_r2_1,
       r2(2) => DANGLING_U5_r2_2,
       r2(3) => DANGLING_U5_r2_3,
       r2(4) => DANGLING_U5_r2_4,
       r2(5) => DANGLING_U5_r2_5,
       r2(6) => DANGLING_U5_r2_6,
       r2(7) => DANGLING_U5_r2_7,
       r2(8) => DANGLING_U5_r2_8,
       r2(9) => DANGLING_U5_r2_9,
       r2(10) => DANGLING_U5_r2_10,
       r2(11) => DANGLING_U5_r2_11,
       r2(12) => DANGLING_U5_r2_12,
       r2(13) => DANGLING_U5_r2_13,
       r2(14) => DANGLING_U5_r2_14,
       r2(15) => DANGLING_U5_r2_15,
       r2(16) => DANGLING_U5_r2_16,
       r2(17) => DANGLING_U5_r2_17,
       r2(18) => DANGLING_U5_r2_18,
       r2(19) => DANGLING_U5_r2_19,
       r2(20) => DANGLING_U5_r2_20,
       r2(21) => DANGLING_U5_r2_21,
       r2(22) => DANGLING_U5_r2_22,
       r2(23) => DANGLING_U5_r2_23,
       r2(24) => DANGLING_U5_r2_24,
       r2(25) => DANGLING_U5_r2_25,
       r2(26) => DANGLING_U5_r2_26,
       r2(27) => DANGLING_U5_r2_27,
       r2(28) => DANGLING_U5_r2_28,
       r2(29) => DANGLING_U5_r2_29,
       r2(30) => DANGLING_U5_r2_30,
       r2(31) => DANGLING_U5_r2_31,
       r2(32) => DANGLING_U5_r2_32,
       r2(33) => DANGLING_U5_r2_33,
       r2(34) => DANGLING_U5_r2_34,
       r2(35) => DANGLING_U5_r2_35,
       r2(36) => DANGLING_U5_r2_36,
       r2(37) => DANGLING_U5_r2_37,
       r2(38) => DANGLING_U5_r2_38,
       r2(39) => DANGLING_U5_r2_39,
       r2(40) => DANGLING_U5_r2_40,
       r2(41) => DANGLING_U5_r2_41,
       r2(42) => DANGLING_U5_r2_42,
       r2(43) => DANGLING_U5_r2_43,
       r2(44) => DANGLING_U5_r2_44,
       r2(45) => DANGLING_U5_r2_45,
       r2(46) => DANGLING_U5_r2_46,
       r2(47) => DANGLING_U5_r2_47,
       r2(48) => DANGLING_U5_r2_48,
       r2(49) => DANGLING_U5_r2_49,
       r2(50) => DANGLING_U5_r2_50,
       r2(51) => DANGLING_U5_r2_51,
       r2(52) => DANGLING_U5_r2_52,
       r2(53) => DANGLING_U5_r2_53,
       r2(54) => DANGLING_U5_r2_54,
       r2(55) => DANGLING_U5_r2_55,
       r2(56) => DANGLING_U5_r2_56,
       r2(57) => DANGLING_U5_r2_57,
       r2(58) => DANGLING_U5_r2_58,
       r2(59) => DANGLING_U5_r2_59,
       r2(60) => DANGLING_U5_r2_60,
       r2(61) => DANGLING_U5_r2_61,
       r2(62) => DANGLING_U5_r2_62,
       r2(63) => DANGLING_U5_r2_63,
       r2(64) => DANGLING_U5_r2_64,
       r2(65) => DANGLING_U5_r2_65,
       r2(66) => DANGLING_U5_r2_66,
       r2(67) => DANGLING_U5_r2_67,
       r2(68) => DANGLING_U5_r2_68,
       r2(69) => DANGLING_U5_r2_69,
       r2(70) => DANGLING_U5_r2_70,
       r2(71) => DANGLING_U5_r2_71,
       r2(72) => DANGLING_U5_r2_72,
       r2(73) => DANGLING_U5_r2_73,
       r2(74) => DANGLING_U5_r2_74,
       r2(75) => DANGLING_U5_r2_75,
       r2(76) => DANGLING_U5_r2_76,
       r2(77) => DANGLING_U5_r2_77,
       r2(78) => DANGLING_U5_r2_78,
       r2(79) => DANGLING_U5_r2_79,
       r2(80) => DANGLING_U5_r2_80,
       r2(81) => DANGLING_U5_r2_81,
       r2(82) => DANGLING_U5_r2_82,
       r2(83) => DANGLING_U5_r2_83,
       r2(84) => DANGLING_U5_r2_84,
       r2(85) => DANGLING_U5_r2_85,
       r2(86) => DANGLING_U5_r2_86,
       r2(87) => DANGLING_U5_r2_87,
       r2(88) => DANGLING_U5_r2_88,
       r2(89) => DANGLING_U5_r2_89,
       r2(90) => DANGLING_U5_r2_90,
       r2(91) => DANGLING_U5_r2_91,
       r2(92) => DANGLING_U5_r2_92,
       r2(93) => DANGLING_U5_r2_93,
       r2(94) => DANGLING_U5_r2_94,
       r2(95) => DANGLING_U5_r2_95,
       r2(96) => DANGLING_U5_r2_96,
       r2(97) => DANGLING_U5_r2_97,
       r2(98) => DANGLING_U5_r2_98,
       r2(99) => DANGLING_U5_r2_99,
       r2(100) => DANGLING_U5_r2_100,
       r2(101) => DANGLING_U5_r2_101,
       r2(102) => DANGLING_U5_r2_102,
       r2(103) => DANGLING_U5_r2_103,
       r2(104) => DANGLING_U5_r2_104,
       r2(105) => DANGLING_U5_r2_105,
       r2(106) => DANGLING_U5_r2_106,
       r2(107) => DANGLING_U5_r2_107,
       r2(108) => DANGLING_U5_r2_108,
       r2(109) => DANGLING_U5_r2_109,
       r2(110) => DANGLING_U5_r2_110,
       r2(111) => DANGLING_U5_r2_111,
       r2(112) => DANGLING_U5_r2_112,
       r2(113) => DANGLING_U5_r2_113,
       r2(114) => DANGLING_U5_r2_114,
       r2(115) => DANGLING_U5_r2_115,
       r2(116) => DANGLING_U5_r2_116,
       r2(117) => DANGLING_U5_r2_117,
       r2(118) => DANGLING_U5_r2_118,
       r2(119) => DANGLING_U5_r2_119,
       r2(120) => DANGLING_U5_r2_120,
       r2(121) => DANGLING_U5_r2_121,
       r2(122) => DANGLING_U5_r2_122,
       r2(123) => DANGLING_U5_r2_123,
       r2(124) => DANGLING_U5_r2_124,
       r2(125) => DANGLING_U5_r2_125,
       r2(126) => DANGLING_U5_r2_126,
       r2(127) => NET134,
       r3(0) => DANGLING_U5_r3_0,
       r3(1) => DANGLING_U5_r3_1,
       r3(2) => DANGLING_U5_r3_2,
       r3(3) => DANGLING_U5_r3_3,
       r3(4) => DANGLING_U5_r3_4,
       r3(5) => DANGLING_U5_r3_5,
       r3(6) => DANGLING_U5_r3_6,
       r3(7) => DANGLING_U5_r3_7,
       r3(8) => DANGLING_U5_r3_8,
       r3(9) => DANGLING_U5_r3_9,
       r3(10) => DANGLING_U5_r3_10,
       r3(11) => DANGLING_U5_r3_11,
       r3(12) => DANGLING_U5_r3_12,
       r3(13) => DANGLING_U5_r3_13,
       r3(14) => DANGLING_U5_r3_14,
       r3(15) => DANGLING_U5_r3_15,
       r3(16) => DANGLING_U5_r3_16,
       r3(17) => DANGLING_U5_r3_17,
       r3(18) => DANGLING_U5_r3_18,
       r3(19) => DANGLING_U5_r3_19,
       r3(20) => DANGLING_U5_r3_20,
       r3(21) => DANGLING_U5_r3_21,
       r3(22) => DANGLING_U5_r3_22,
       r3(23) => DANGLING_U5_r3_23,
       r3(24) => DANGLING_U5_r3_24,
       r3(25) => DANGLING_U5_r3_25,
       r3(26) => DANGLING_U5_r3_26,
       r3(27) => DANGLING_U5_r3_27,
       r3(28) => DANGLING_U5_r3_28,
       r3(29) => DANGLING_U5_r3_29,
       r3(30) => DANGLING_U5_r3_30,
       r3(31) => DANGLING_U5_r3_31,
       r3(32) => DANGLING_U5_r3_32,
       r3(33) => DANGLING_U5_r3_33,
       r3(34) => DANGLING_U5_r3_34,
       r3(35) => DANGLING_U5_r3_35,
       r3(36) => DANGLING_U5_r3_36,
       r3(37) => DANGLING_U5_r3_37,
       r3(38) => DANGLING_U5_r3_38,
       r3(39) => DANGLING_U5_r3_39,
       r3(40) => DANGLING_U5_r3_40,
       r3(41) => DANGLING_U5_r3_41,
       r3(42) => DANGLING_U5_r3_42,
       r3(43) => DANGLING_U5_r3_43,
       r3(44) => DANGLING_U5_r3_44,
       r3(45) => DANGLING_U5_r3_45,
       r3(46) => DANGLING_U5_r3_46,
       r3(47) => DANGLING_U5_r3_47,
       r3(48) => DANGLING_U5_r3_48,
       r3(49) => DANGLING_U5_r3_49,
       r3(50) => DANGLING_U5_r3_50,
       r3(51) => DANGLING_U5_r3_51,
       r3(52) => DANGLING_U5_r3_52,
       r3(53) => DANGLING_U5_r3_53,
       r3(54) => DANGLING_U5_r3_54,
       r3(55) => DANGLING_U5_r3_55,
       r3(56) => DANGLING_U5_r3_56,
       r3(57) => DANGLING_U5_r3_57,
       r3(58) => DANGLING_U5_r3_58,
       r3(59) => DANGLING_U5_r3_59,
       r3(60) => DANGLING_U5_r3_60,
       r3(61) => DANGLING_U5_r3_61,
       r3(62) => DANGLING_U5_r3_62,
       r3(63) => DANGLING_U5_r3_63,
       r3(64) => DANGLING_U5_r3_64,
       r3(65) => DANGLING_U5_r3_65,
       r3(66) => DANGLING_U5_r3_66,
       r3(67) => DANGLING_U5_r3_67,
       r3(68) => DANGLING_U5_r3_68,
       r3(69) => DANGLING_U5_r3_69,
       r3(70) => DANGLING_U5_r3_70,
       r3(71) => DANGLING_U5_r3_71,
       r3(72) => DANGLING_U5_r3_72,
       r3(73) => DANGLING_U5_r3_73,
       r3(74) => DANGLING_U5_r3_74,
       r3(75) => DANGLING_U5_r3_75,
       r3(76) => DANGLING_U5_r3_76,
       r3(77) => DANGLING_U5_r3_77,
       r3(78) => DANGLING_U5_r3_78,
       r3(79) => DANGLING_U5_r3_79,
       r3(80) => DANGLING_U5_r3_80,
       r3(81) => DANGLING_U5_r3_81,
       r3(82) => DANGLING_U5_r3_82,
       r3(83) => DANGLING_U5_r3_83,
       r3(84) => DANGLING_U5_r3_84,
       r3(85) => DANGLING_U5_r3_85,
       r3(86) => DANGLING_U5_r3_86,
       r3(87) => DANGLING_U5_r3_87,
       r3(88) => DANGLING_U5_r3_88,
       r3(89) => DANGLING_U5_r3_89,
       r3(90) => DANGLING_U5_r3_90,
       r3(91) => DANGLING_U5_r3_91,
       r3(92) => DANGLING_U5_r3_92,
       r3(93) => DANGLING_U5_r3_93,
       r3(94) => DANGLING_U5_r3_94,
       r3(95) => DANGLING_U5_r3_95,
       r3(96) => DANGLING_U5_r3_96,
       r3(97) => DANGLING_U5_r3_97,
       r3(98) => DANGLING_U5_r3_98,
       r3(99) => DANGLING_U5_r3_99,
       r3(100) => DANGLING_U5_r3_100,
       r3(101) => DANGLING_U5_r3_101,
       r3(102) => DANGLING_U5_r3_102,
       r3(103) => DANGLING_U5_r3_103,
       r3(104) => DANGLING_U5_r3_104,
       r3(105) => DANGLING_U5_r3_105,
       r3(106) => DANGLING_U5_r3_106,
       r3(107) => DANGLING_U5_r3_107,
       r3(108) => DANGLING_U5_r3_108,
       r3(109) => DANGLING_U5_r3_109,
       r3(110) => DANGLING_U5_r3_110,
       r3(111) => DANGLING_U5_r3_111,
       r3(112) => DANGLING_U5_r3_112,
       r3(113) => DANGLING_U5_r3_113,
       r3(114) => DANGLING_U5_r3_114,
       r3(115) => DANGLING_U5_r3_115,
       r3(116) => DANGLING_U5_r3_116,
       r3(117) => DANGLING_U5_r3_117,
       r3(118) => DANGLING_U5_r3_118,
       r3(119) => DANGLING_U5_r3_119,
       r3(120) => DANGLING_U5_r3_120,
       r3(121) => DANGLING_U5_r3_121,
       r3(122) => DANGLING_U5_r3_122,
       r3(123) => DANGLING_U5_r3_123,
       r3(124) => DANGLING_U5_r3_124,
       r3(125) => DANGLING_U5_r3_125,
       r3(126) => DANGLING_U5_r3_126,
       r3(127) => NET168,
       WrData(0) => Dangling_Input_Signal,
       WrData(1) => Dangling_Input_Signal,
       WrData(2) => Dangling_Input_Signal,
       WrData(3) => Dangling_Input_Signal,
       WrData(4) => Dangling_Input_Signal,
       WrData(5) => Dangling_Input_Signal,
       WrData(6) => Dangling_Input_Signal,
       WrData(7) => Dangling_Input_Signal,
       WrData(8) => Dangling_Input_Signal,
       WrData(9) => Dangling_Input_Signal,
       WrData(10) => Dangling_Input_Signal,
       WrData(11) => Dangling_Input_Signal,
       WrData(12) => Dangling_Input_Signal,
       WrData(13) => Dangling_Input_Signal,
       WrData(14) => Dangling_Input_Signal,
       WrData(15) => Dangling_Input_Signal,
       WrData(16) => Dangling_Input_Signal,
       WrData(17) => Dangling_Input_Signal,
       WrData(18) => Dangling_Input_Signal,
       WrData(19) => Dangling_Input_Signal,
       WrData(20) => Dangling_Input_Signal,
       WrData(21) => Dangling_Input_Signal,
       WrData(22) => Dangling_Input_Signal,
       WrData(23) => Dangling_Input_Signal,
       WrData(24) => Dangling_Input_Signal,
       WrData(25) => Dangling_Input_Signal,
       WrData(26) => Dangling_Input_Signal,
       WrData(27) => Dangling_Input_Signal,
       WrData(28) => Dangling_Input_Signal,
       WrData(29) => Dangling_Input_Signal,
       WrData(30) => Dangling_Input_Signal,
       WrData(31) => Dangling_Input_Signal,
       WrData(32) => Dangling_Input_Signal,
       WrData(33) => Dangling_Input_Signal,
       WrData(34) => Dangling_Input_Signal,
       WrData(35) => Dangling_Input_Signal,
       WrData(36) => Dangling_Input_Signal,
       WrData(37) => Dangling_Input_Signal,
       WrData(38) => Dangling_Input_Signal,
       WrData(39) => Dangling_Input_Signal,
       WrData(40) => Dangling_Input_Signal,
       WrData(41) => Dangling_Input_Signal,
       WrData(42) => Dangling_Input_Signal,
       WrData(43) => Dangling_Input_Signal,
       WrData(44) => Dangling_Input_Signal,
       WrData(45) => Dangling_Input_Signal,
       WrData(46) => Dangling_Input_Signal,
       WrData(47) => Dangling_Input_Signal,
       WrData(48) => Dangling_Input_Signal,
       WrData(49) => Dangling_Input_Signal,
       WrData(50) => Dangling_Input_Signal,
       WrData(51) => Dangling_Input_Signal,
       WrData(52) => Dangling_Input_Signal,
       WrData(53) => Dangling_Input_Signal,
       WrData(54) => Dangling_Input_Signal,
       WrData(55) => Dangling_Input_Signal,
       WrData(56) => Dangling_Input_Signal,
       WrData(57) => Dangling_Input_Signal,
       WrData(58) => Dangling_Input_Signal,
       WrData(59) => Dangling_Input_Signal,
       WrData(60) => Dangling_Input_Signal,
       WrData(61) => Dangling_Input_Signal,
       WrData(62) => Dangling_Input_Signal,
       WrData(63) => Dangling_Input_Signal,
       WrData(64) => Dangling_Input_Signal,
       WrData(65) => Dangling_Input_Signal,
       WrData(66) => Dangling_Input_Signal,
       WrData(67) => Dangling_Input_Signal,
       WrData(68) => Dangling_Input_Signal,
       WrData(69) => Dangling_Input_Signal,
       WrData(70) => Dangling_Input_Signal,
       WrData(71) => Dangling_Input_Signal,
       WrData(72) => Dangling_Input_Signal,
       WrData(73) => Dangling_Input_Signal,
       WrData(74) => Dangling_Input_Signal,
       WrData(75) => Dangling_Input_Signal,
       WrData(76) => Dangling_Input_Signal,
       WrData(77) => Dangling_Input_Signal,
       WrData(78) => Dangling_Input_Signal,
       WrData(79) => Dangling_Input_Signal,
       WrData(80) => Dangling_Input_Signal,
       WrData(81) => Dangling_Input_Signal,
       WrData(82) => Dangling_Input_Signal,
       WrData(83) => Dangling_Input_Signal,
       WrData(84) => Dangling_Input_Signal,
       WrData(85) => Dangling_Input_Signal,
       WrData(86) => Dangling_Input_Signal,
       WrData(87) => Dangling_Input_Signal,
       WrData(88) => Dangling_Input_Signal,
       WrData(89) => Dangling_Input_Signal,
       WrData(90) => Dangling_Input_Signal,
       WrData(91) => Dangling_Input_Signal,
       WrData(92) => Dangling_Input_Signal,
       WrData(93) => Dangling_Input_Signal,
       WrData(94) => Dangling_Input_Signal,
       WrData(95) => Dangling_Input_Signal,
       WrData(96) => Dangling_Input_Signal,
       WrData(97) => Dangling_Input_Signal,
       WrData(98) => Dangling_Input_Signal,
       WrData(99) => Dangling_Input_Signal,
       WrData(100) => Dangling_Input_Signal,
       WrData(101) => Dangling_Input_Signal,
       WrData(102) => Dangling_Input_Signal,
       WrData(103) => Dangling_Input_Signal,
       WrData(104) => Dangling_Input_Signal,
       WrData(105) => Dangling_Input_Signal,
       WrData(106) => Dangling_Input_Signal,
       WrData(107) => Dangling_Input_Signal,
       WrData(108) => Dangling_Input_Signal,
       WrData(109) => Dangling_Input_Signal,
       WrData(110) => Dangling_Input_Signal,
       WrData(111) => Dangling_Input_Signal,
       WrData(112) => Dangling_Input_Signal,
       WrData(113) => Dangling_Input_Signal,
       WrData(114) => Dangling_Input_Signal,
       WrData(115) => Dangling_Input_Signal,
       WrData(116) => Dangling_Input_Signal,
       WrData(117) => Dangling_Input_Signal,
       WrData(118) => Dangling_Input_Signal,
       WrData(119) => Dangling_Input_Signal,
       WrData(120) => Dangling_Input_Signal,
       WrData(121) => Dangling_Input_Signal,
       WrData(122) => Dangling_Input_Signal,
       WrData(123) => Dangling_Input_Signal,
       WrData(124) => Dangling_Input_Signal,
       WrData(125) => Dangling_Input_Signal,
       WrData(126) => Dangling_Input_Signal,
       WrData(127) => NET210,
       clk => clk
  );


---- Dangling input signal assignment ----

Dangling_Input_Signal <= DANGLING_INPUT_CONSTANT;

end block_diagram;
